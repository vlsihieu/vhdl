----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    01:39:34 12/04/2019 
-- Design Name: 
-- Module Name:    LCD_20X4_GAN_DULIEU_1SO_TO - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LCD_20X4_GAN_DULIEU_1SO_TO is
    Port ( 
			  lcd_so_X   : in  STD_LOGIC_VECTOR (47 downto 0);
			  -----------------------------------------
			  H2_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  H2_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  H1_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  H1_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  H1_18 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  H1_19 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			  -----------------------------------------
			  ena_8led : in std_logic_vector(7 downto 0);
			  ena_4led : in std_logic_vector(3 downto 0);
			  -------------------------------------------
			  ena1hz : in std_logic;
			  rst    : in std_logic;
			  --------------------------------------------
           LCD_H1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H2 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H3 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H4 : out  STD_LOGIC_VECTOR (159 downto 0));
end LCD_20X4_GAN_DULIEU_1SO_TO;

architecture Behavioral of LCD_20X4_GAN_DULIEU_1SO_TO is
TYPE MANG_DICH IS ARRAY(INTEGER RANGE 0 TO 25) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL HOVATEN : MANG_DICH:= ( 

      0  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8), 
		1  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		2  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		3  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		4  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		5  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		6  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		7  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		8  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		9  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
---------------------------------------      
      13  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8), 
      14  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),
	   15  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8),
	   16  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8),
		17  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		18  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8),
		19  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),
		20  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8),
		21  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		22  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('B'),8),
		23  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8),
		24  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8),
		25  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8)
		);
begin
	 PROCESS(RST,ENA1hz,HOVATEN)
	 BEGIN
		IF (RST = '1') THEN 	HOVATEN <=(
      0  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8), 
		1  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		2  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		3  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		4  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		5  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		6  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		7  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		8  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		9  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		10 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		11 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		12 => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
---------------------------------------      
      13  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8), 
      14  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8),
	   15  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8),
	   16  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8),
		17  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		18  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8),
		19  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8),
		20  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8),
		21  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8),
		22  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('B'),8),
		23  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8),
		24  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8),
		25  => CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8)
      );
		ELSIF (FALLING_EDGE(ENA1HZ)) THEN
			HOVATEN(25) <= HOVATEN(0);
			FOR I IN 0 TO 24
			LOOP
				HOVATEN(I) <= HOVATEN(I+1);
			END LOOP;
		ELSE
			HOVATEN <= HOVATEN;
		END IF;
	 END PROCESS;


---- HANG 1
	LCD_H1(  7 DOWNTO   0) 		<= X"3" & H1_0 when ena_4led(0) = '1' else
	                              X"20";
	LCD_H1( 15 DOWNTO   8) 		<= X"3" & H1_1 WHEN ena_4led(1) = '1' else
	                              X"20";
	LCD_H1( 23 DOWNTO  16) 		<= lcd_so_X (47 DOWNTO 40);
	LCD_H1( 31 DOWNTO  24) 		<= lcd_so_X (39 DOWNTO 32);
	LCD_H1( 39 DOWNTO  32) 		<= lcd_so_X (31 DOWNTO 24);
	LCD_H1( 47 DOWNTO  40) 		<= HOVATEN(0);
	LCD_H1( 55 DOWNTO  48) 		<= HOVATEN(1);
	LCD_H1( 63 DOWNTO  56) 		<= HOVATEN(2);
	LCD_H1( 71 DOWNTO  64) 		<= HOVATEN(3);
	LCD_H1( 79 DOWNTO  72) 		<= HOVATEN(4);
	LCD_H1( 87 DOWNTO  80) 		<= HOVATEN(5);
	LCD_H1( 95 DOWNTO  88) 		<= HOVATEN(6);
	LCD_H1(103 DOWNTO  96) 		<= HOVATEN(7);
	LCD_H1(111 DOWNTO 104) 		<= HOVATEN(8);
	LCD_H1(119 DOWNTO 112) 		<= HOVATEN(9);
	LCD_H1(127 DOWNTO 120) 		<= HOVATEN(10);
	LCD_H1(135 DOWNTO 128) 		<= HOVATEN(11);
	LCD_H1(143 DOWNTO 136) 		<= HOVATEN(12);
	LCD_H1(151 DOWNTO 144) 		<= X"3" & H1_18;
	LCD_H1(159 DOWNTO 152) 		<= X"3" & H1_19;
	
---- HANG 2
	LCD_H2(  7 DOWNTO   0) 		<= X"3" & H2_0 WHEN ENA_4LED(2) = '1' ELSE
	                              X"20";
	LCD_H2( 15 DOWNTO   8) 		<= X"3" & H2_1 WHEN ENA_4LED(3) = '1' ELSE
	                              X"20";
	LCD_H2( 23 DOWNTO  16) 		<= lcd_so_X (23 DOWNTO 16);
	LCD_H2( 31 DOWNTO  24) 		<= lcd_so_X (15 DOWNTO 8);
	LCD_H2( 39 DOWNTO  32) 		<= lcd_so_X (7 DOWNTO 0);
	LCD_H2( 47 DOWNTO  40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8) WHEN ena_8led(7) ='1' else
	                              X"20";
	LCD_H2( 55 DOWNTO  48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('6'),8) WHEN ENA_8LED(6) = '1' ELSE
	                              X"20";
	LCD_H2( 63 DOWNTO  56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8) WHEN ENA_8LED(5) = '1' ELSE
	                              X"20";
	LCD_H2( 71 DOWNTO  64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8) WHEN ENA_8LED(4) = '1' ELSE
	                              X"20";
	LCD_H2( 79 DOWNTO  72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('9'),8) WHEN ENA_8LED(3) = '1' ELSE
	                              X"20";
	LCD_H2( 87 DOWNTO  80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('0'),8) WHEN ENA_8LED(2) = '1' ELSE
	                              X"20";
	LCD_H2( 95 DOWNTO  88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('8'),8) WHEN ENA_8LED(1) = '1' ELSE
	                              X"20";
	LCD_H2(103 DOWNTO  96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('8'),8) WHEN ENA_8LED(0) = '1' ELSE
	                              X"20";
	LCD_H2(111 DOWNTO 104) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(119 DOWNTO 112) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(127 DOWNTO 120) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(135 DOWNTO 128) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(143 DOWNTO 136) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(151 DOWNTO 144) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(159 DOWNTO 152) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	
---- HANG 3
	LCD_H3(  7 DOWNTO   0) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_H3( 15 DOWNTO   8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_H3( 23 DOWNTO  16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	LCD_H3( 31 DOWNTO  24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3( 39 DOWNTO  32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_H3( 47 DOWNTO  40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_H3( 55 DOWNTO  48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_H3( 63 DOWNTO  56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3( 71 DOWNTO  64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('S'),8);
	LCD_H3( 79 DOWNTO  72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('P'),8);
	LCD_H3( 87 DOWNTO  80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_H3( 95 DOWNTO  88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_H3(103 DOWNTO  96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3(111 DOWNTO 104) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_H3(119 DOWNTO 112) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_H3(127 DOWNTO 120) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_H3(135 DOWNTO 128) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_H3(143 DOWNTO 136) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('5'),8);
	LCD_H3(151 DOWNTO 144) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('6'),8);
	LCD_H3(159 DOWNTO 152) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('7'),8);
	
---- HANG 4
	LCD_H4(  7 DOWNTO   0) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_H4( 15 DOWNTO   8) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_H4( 23 DOWNTO  16) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	LCD_H4( 31 DOWNTO  24) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4( 39 DOWNTO  32) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_H4( 47 DOWNTO  40) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_H4( 55 DOWNTO  48) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_H4( 63 DOWNTO  56) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4( 71 DOWNTO  64) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('S'),8);
	LCD_H4( 79 DOWNTO  72) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('P'),8);
	LCD_H4( 87 DOWNTO  80) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_H4( 95 DOWNTO  88) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_H4(103 DOWNTO  96) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(111 DOWNTO 104) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('7'),8);
	LCD_H4(119 DOWNTO 112) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('6'),8);
	LCD_H4(127 DOWNTO 120) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('5'),8);
	LCD_H4(135 DOWNTO 128) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_H4(143 DOWNTO 136) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_H4(151 DOWNTO 144) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_H4(159 DOWNTO 152) 		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);



end Behavioral;

