library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;



entity DIEUKHIEN_MODE is
	 Port ( SEL_3B : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
           RST: IN STD_LOGIC;
           OE : out  STD_LOGIC_VECTOR(3 DOWNTO 0)
			  );
end DIEUKHIEN_MODE;

architecture Behavioral of DIEUKHIEN_MODE is
begin
	PROCESS(SEL_3B,RST)
	BEGIN
	   OE <= "0000";
		IF RST = '1' THEN OE <= "0000";
		ELSIF (SEL_3B = "000") THEN OE <="0000";
		ELSIF (SEL_3B = "001") THEN OE <="0001";
		ELSIF (SEL_3B = "010") THEN OE <="0010";
		ELSIF (SEL_3B = "011") THEN OE <="0100";
		ELSIF (SEL_3B = "100") THEN OE <="1000";
		END IF;
	END PROCESS;

end Behavioral;