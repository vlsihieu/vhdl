-- CHUONG TRINH CHIA XUNG CHO CAC BAI

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CHIA_10ENA IS 
	PORT( CKHT: IN STD_LOGIC;
			OE : IN STD_LOGIC_VECTOR( 1 DOWNTO 0 );
			ENA_CK : OUT STD_LOGIC);
END CHIA_10ENA;
 
ARCHITECTURE BEHAVIORAL OF CHIA_10ENA IS

--SIGNAL ENA2HZ  : STD_LOGIC; 
SIGNAL ENA5HZ  : STD_LOGIC;  
SIGNAL ENA10HZ  : STD_LOGIC; 

CONSTANT N : INTEGER := 50000000;


SIGNAL D10HZ_REG,  D10HZ_NEXT  : INTEGER RANGE 0 TO N/10 := 1;
SIGNAL D5HZ_REG,   D5HZ_NEXT   : INTEGER RANGE 0 TO N/5 := 1;
--SIGNAL D2HZ_REG,   D2HZ_NEXT   : INTEGER RANGE 0 TO N/2 := 1;

BEGIN
-- OUTPUT LOGIC

--	ENA2HZ   <='1' WHEN D2HZ_REG = N/(2*2)  	  	ELSE '0';
	ENA5HZ   <='1' WHEN D5HZ_REG = N/(5*2)        ELSE '0';
	ENA10HZ  <='1' WHEN D10HZ_REG = N/(10*2)      ELSE '0';  


	
-- REGISTER
PROCESS( CKHT)
BEGIN	
		IF FALLING_EDGE (CKHT) THEN D10HZ_REG   <= D10HZ_NEXT;
											 D5HZ_REG    <= D5HZ_NEXT;
--											 D2HZ_REG    <= D2HZ_NEXT;

		END IF;
	END PROCESS;
	
-- NEXT STATE LOGIC

						


D10HZ_NEXT <= 1 WHEN D10HZ_REG = N/10 ELSE
						D10HZ_REG +1;  

D5HZ_NEXT <= 1 WHEN D5HZ_REG = N/5 ELSE
						D5HZ_REG +1;
--
--D2HZ_NEXT <= 1 WHEN D2HZ_REG = N/2 ELSE
--						D2HZ_REG +1;


-- PHAN CHIA XUNG CHO TUNG BAI 

ENA_CK <= ENA10HZ WHEN OE = "01" ELSE	-- PST 10HZ
			 ENA5HZ  WHEN OE = "10" ELSE  -- TSP 5HZ
--			 ENA2HZ  WHEN OE = "100" ELSE  -- DS 1 LED 2HZ
			 '0' ;
			
						
	
END BEHAVIORAL;
	