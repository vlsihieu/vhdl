library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
entity XULY_MOD is
    Port ( CKHT, ENA_DB: in  STD_LOGIC;
           GIATRI_MOD: OUT  STD_LOGIC_VECTOR(1 DOWNTO 0)
			  );
end XULY_MOD;

architecture Behavioral of XULY_MOD is
SIGNAL GIATRI_MOD_REG:  STD_LOGIC_VECTOR(1 DOWNTO 0):="00";
SIGNAL GIATRI_MOD_NEXT:  STD_LOGIC_VECTOR(1 DOWNTO 0);
begin
	PROCESS (CKHT)
   BEGIN   
       IF FALLING_EDGE(CKHT) THEN GIATRI_MOD_REG <= GIATRI_MOD_NEXT;
		 END IF;
	END PROCESS;
		 
	GIATRI_MOD_NEXT <= 	GIATRI_MOD_REG + 1 WHEN ENA_DB = '1' ELSE
								GIATRI_MOD_REG;
	 
	GIATRI_MOD <= GIATRI_MOD_REG;
end Behavioral;