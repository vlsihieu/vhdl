LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;



ENTITY LED_STD_TNV_TTR IS
PORT ( CKHT : IN STD_LOGIC;
       RST : IN STD_LOGIC;
		 ENA_DB  :IN STD_LOGIC;
		 ENA_SS: IN STD_LOGIC;
		 DEM: IN STD_LOGIC;
		 Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END LED_STD_TNV_TTR;

ARCHITECTURE THAN OF LED_STD_TNV_TTR IS
SIGNAL Q_R, Q_N: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN Q_R <= (OTHERS => '0');
	ELSIF FALLING_EDGE(CKHT) THEN Q_R<=Q_N;
	END IF;
END PROCESS;

PROCESS(ENA_DB,DEM,ENA_SS,Q_R)
BEGIN
	Q_N <= Q_R;
	IF ENA_DB = '1' THEN
	  IF ENA_SS = '1' THEN 
		 IF DEM = '0' THEN 
             Q_N<= NOT(Q_R(4)) & Q_R(7 DOWNTO 5) & Q_R(2 DOWNTO 0) & NOT(Q_R(3));
		 ELSIF DEM = '1' THEN 
			    Q_N<= Q_R(6 DOWNTO 4) & NOT(Q_R(7)) & NOT(Q_R(0)) & Q_R(3 DOWNTO 1);
		 END IF;
	  END IF;
	END IF;
END PROCESS;
	Q <= Q_R;		
--Q <= Q_REG WHEN ENA_SS = '1' ELSE (OTHERS => '0');
END THAN;
