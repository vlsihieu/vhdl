LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY MACHDEM_GH IS 
	PORT (     CKHT,RST : IN STD_LOGIC;
				  ENA_DB   : IN STd_LOGIC;
				  GH_DV_TREN: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
				  GH_DV_DUOI: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
				  GH_CHUC_TREN: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
				  GH_CHUC_DUOI : IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
				  DONVI,CHUC: OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0));
END MACHDEM_GH;
ARCHITECTURE PMH OF MACHDEM_GH IS 
SIGNAL DONVI_REG:STD_LOGIC_VECTOR(3 DOWNTO 0) := GH_DV_DUOI;
signal DONVI_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG :STD_LOGIC_VECTOR(3 DOWNTO 0):= GH_CHUC_DUOI;
signal CHUC_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0 );
BEGIN
	PROCESS (CKHT, RST,GH_DV_DUOI,GH_CHUC_DUOI)
	BEGIN
		IF RST='1' THEN DONVI_REG <= GH_DV_DUOI;			
							 CHUC_REG <= GH_CHUC_DUOI;
		ELSIF FALLING_EDGE (CKHT) THEN DONVI_REG <= DONVI_NEXT;
												 CHUC_REG <= CHUC_NEXT;
		END IF;
	END PROCESS;
	PROCESS (DONVI_REG, CHUC_REG,  ENA_DB ,GH_DV_DUOI,GH_DV_TREN,GH_CHUC_DUOI,GH_CHUC_TREN)
	BEGIN
		DONVI_NEXT <= DONVI_REG;
		CHUC_NEXT <= CHUC_REG;
		IF ENA_DB ='1' THEN 
			IF (GH_CHUC_TREN < GH_CHUC_DUOI )  or (gh_dv_tren < gh_dv_duoi) THEN DONVI_NEXT <= GH_DV_DUOI;	
													                   CHUC_NEXT  <= GH_CHUC_DUOI;
			ELSif (GH_CHUC_TREN > GH_CHUC_DUOI) or (gh_dv_tren > gh_dv_duoi) then
				IF DONVI_REG = GH_DV_TREN AND CHUC_REG = GH_CHUC_TREN THEN DONVI_NEXT <= GH_DV_DUOI;
																							  CHUC_NEXT  <= GH_CHUC_DUOI;
				ELSE 																		
					IF DONVI_REG /= X"9" THEN DONVI_NEXT <= DONVI_REG +1;
					ELSE							  DONVI_NEXT <= X"0";
						IF CHUC_REG /= X"9" THEN CHUC_NEXT <= CHUC_REG +1;
						ELSE 							 CHUC_NEXT <= X"0";
						END IF;
					END IF;
				END IF;
			END IF;
		END IF;
	END PROCESS;	
	DONVI <= DONVI_REG;
	CHUC <= CHUC_REG;
END PMH;