LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY BTN IS
	PORT ( CKHT: IN STD_LOGIC;
			 BTN: IN STD_LOGIC;
			 Q: OUT STD_LOGIC
		   );
END BTN;

ARCHITECTURE BEHAVIOR OF BTN IS
CONSTANT N: INTEGER:=20;
TYPE DB_STATE IS (ZERO,WAIT0,ONE,WAIT1);
SIGNAL DB_REG,DB_NEXT : DB_STATE;

SIGNAL QFF,DB_TICK : STD_LOGIC;
SIGNAL DELAY_REG, DELAY_NEXT: UNSIGNED (N-1 DOWNTO 0);
BEGIN
PROCESS (CKHT)
BEGIN
	IF FALLING_EDGE (CKHT) THEN DB_REG <= DB_NEXT;
										 DELAY_REG <= DELAY_NEXT;
										 QFF <= DB_TICK;
	END IF;
END PROCESS;
PROCESS(DELAY_REG,DELAY_NEXT,BTN)
BEGIN
	DELAY_NEXT <= DELAY_REG;
	DB_NEXT <= DB_REG;
	CASE DB_REG IS
		WHEN ZERO => DB_TICK <= '0';
						 IF (BTN = '1') THEN DB_NEXT <= WAIT1;
												  DELAY_NEXT <= (OTHERS => '1');
						 END IF;
		WHEN WAIT1 => DB_TICK <= '0';
						 IF (BTN= '1') THEN DELAY_NEXT <= DELAY_REG -1;
								IF (DELAY_REG =0) THEN DB_NEXT <=ONE;
								END IF;
						 ELSE               DB_NEXT <=ZERO;
						 END IF;
		WHEN ONE => DB_TICK <= '1';
						 IF (BTN= '0') THEN DB_NEXT <= WAIT0;
												  DELAY_NEXT <= (OTHERS => '1');
						 END IF;
		WHEN WAIT0 => DB_TICK <= '1';
						 IF (BTN= '0') THEN DELAY_NEXT <= DELAY_REG -1;
								IF (DELAY_REG =0) THEN DB_NEXT <=ZERO;
								END IF;
						 ELSE               DB_NEXT <=ONE;
						 END IF;	
      END CASE;					 
END PROCESS;
Q <= (NOT QFF) AND DB_TICK;
-- q <= db_tick;
END BEHAVIOR;