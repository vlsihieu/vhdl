library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LCD_20X4_GAN_DULIEU_1SO_TO is
    Port ( ENA_TN:IN STD_LOGIC;
			  H1_19 : in  STD_LOGIC_VECTOR (3 downto 0);
           H1_18 : in  STD_LOGIC_VECTOR (3 downto 0);
           H1_16 : in  STD_LOGIC_VECTOR (3 downto 0);
			  H1_15 : in  STD_LOGIC_VECTOR (3 downto 0);
           H1_13 : in  STD_LOGIC_VECTOR (3 downto 0);
           H1_12 : in  STD_LOGIC_VECTOR (3 downto 0);
			  ND_TRAM,ND_CHUC,ND_DV: IN STD_LOGIC_VECTOR (3 downto 0);
			  LCD_MA_DV_GIO: IN STD_LOGIC_VECTOR(47 DOWNTO 0);
			  LCD_MA_CH_GIO:IN STD_LOGIC_VECTOR(47 DOWNTO 0);
				ENA_CP: IN STD_LOGIC;
			  
			  LCD_MA_TRAM:IN STD_LOGIC_VECTOR(47 DOWNTO 0);
			  LCD_MA_CHUC:IN 	STD_LOGIC_VECTOR(47 DOWNTO 0);
			  LCD_MA_DONVI: IN	STD_LOGIC_VECTOR(47 DOWNTO 0);
           LCD_H1 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H2 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H3 : out  STD_LOGIC_VECTOR (159 downto 0);
           LCD_H4 : out  STD_LOGIC_VECTOR (159 downto 0));
			  
end LCD_20X4_GAN_DULIEU_1SO_TO;

architecture Behavioral of LCD_20X4_GAN_DULIEU_1SO_TO is

begin

--HANG 1
	LCD_H1(7 	DOWNTO 0) 	<= X"20" ;
	LCD_H1(15 	DOWNTO 8) 	<= X"20" ;
	LCD_H1(23	DOWNTO 16) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(47 DOWNTO 40);
	LCD_H1(31 	DOWNTO 24) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(39 DOWNTO 32);
	LCD_H1(39 	DOWNTO 32) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(31 DOWNTO 24);
	LCD_H1(47	DOWNTO 40) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(47 DOWNTO 40);
	LCD_H1(55	DOWNTO 48) 	<= X"3" & H1_12 WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(39 DOWNTO 32);
	LCD_H1(63	DOWNTO 56) 	<= X"3" & H1_13 WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(31 DOWNTO 24);
	LCD_H1(71	DOWNTO 64) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8); 
	LCD_H1(79 	DOWNTO 72) 	<= X"3" & H1_15 ;
	LCD_H1(87 	DOWNTO 80) 	<= X"3" & H1_16 ;
	LCD_H1(95 	DOWNTO 88) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_H1(103 	DOWNTO 96) 	<= X"3" & H1_18 ;
	LCD_H1(111 	DOWNTO 104) <= X"3" & H1_19 ;
	LCD_H1(119	DOWNTO 112) 	<= X"20" ;
	LCD_H1(127 	DOWNTO 120) 	<= X"20";
	LCD_H1(135 	DOWNTO 128) 	<= X"20" ;
	LCD_H1(143	DOWNTO 136) 	<= X"20";
	LCD_H1(151	DOWNTO 144) 	<= X"20" ;
	LCD_H1(159	DOWNTO 152) 	<= X"20" ;

--HANG 2
	LCD_H2(7 	DOWNTO 0) 	<= X"20";
	LCD_H2(15 	DOWNTO 8) 	<= X"20" ;
	LCD_H2(23 	DOWNTO 16) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(23 DOWNTO 16);
	LCD_H2(31 	DOWNTO 24) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(15 DOWNTO 8);
	LCD_H2(39 	DOWNTO 32) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_CH_GIO(7 DOWNTO 0);
	LCD_H2(47	DOWNTO 40) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(23 DOWNTO 16);
	LCD_H2(55 	DOWNTO 48) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(15 DOWNTO 8);
	LCD_H2(63	DOWNTO 56) 	<= X"20" WHEN ENA_TN='0' ELSE LCD_MA_DV_GIO(7 DOWNTO 0);
	LCD_H2(71	DOWNTO 64) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(79 	DOWNTO 72) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(87 	DOWNTO 80) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(95 	DOWNTO 88) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(103 	DOWNTO 96) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(111 	DOWNTO 104) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(119	DOWNTO 112) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(127 	DOWNTO 120) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(135 	DOWNTO 128) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(143	DOWNTO 136) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(151	DOWNTO 144) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H2(159	DOWNTO 152) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	
-- HANG 3
	LCD_H3(7		DOWNTO 0) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_H3(15	DOWNTO 8) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_H3(23	DOWNTO 16) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('I'),8);
	LCD_H3(31	DOWNTO 24) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	LCD_H3(39	DOWNTO 32) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_H3(47	DOWNTO 40) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3(55	DOWNTO 48) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_H3(63	DOWNTO 56) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_H3(71	DOWNTO 64) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3(79	DOWNTO 72) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_H3(87	DOWNTO 80) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H3(95	DOWNTO 88) 	<= X"3" & ND_TRAM WHEN ENA_CP='0' ELSE LCD_MA_TRAM(47 DOWNTO 40);
	LCD_H3(103 	DOWNTO 96) 	<= X"3" & ND_CHUC WHEN ENA_CP='0' ELSE LCD_MA_TRAM(39 DOWNTO 32);
	LCD_H3(111 	DOWNTO 104) <= X"3" & ND_DV   WHEN ENA_CP='0' ELSE LCD_MA_TRAM(31 DOWNTO 24);
										 
	LCD_H3(119 	DOWNTO 112) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(47 DOWNTO 40);
	LCD_H3(127 	DOWNTO 120) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(39 DOWNTO 32);
	LCD_H3(135 	DOWNTO 128) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(31 DOWNTO 24);
									 
	LCD_H3(143 	DOWNTO 136) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_DONVI(47 DOWNTO 40);
	LCD_H3(151 	DOWNTO 144) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_DONVI(39 DOWNTO 32);
	LCD_H3(159 	DOWNTO 152) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_DONVI(31 DOWNTO 24);
	
--HANG 2
	LCD_H4(7 	DOWNTO 0) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(15 	DOWNTO 8) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(23 	DOWNTO 16) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(31	DOWNTO 24) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(39	DOWNTO 32) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(47	DOWNTO 40) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(55	DOWNTO 48) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(63	DOWNTO 56) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(71	DOWNTO 64) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(79 	DOWNTO 72) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(87 	DOWNTO 80) 	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_H4(95	DOWNTO 88) 	<= X"20" WHEN ENA_CP='0' ELSE LCD_MA_TRAM(23 DOWNTO 16);
										
	LCD_H4(103 	DOWNTO 96) 	<= X"20" WHEN ENA_CP='0' ELSE LCD_MA_TRAM(15 DOWNTO 8);
									
	LCD_H4(111 	DOWNTO 104) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_TRAM(7 DOWNTO 0);
									
										 
	LCD_H4(119 	DOWNTO 112) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(23 DOWNTO 16);
	LCD_H4(127 	DOWNTO 120) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(15 DOWNTO 8);
	LCD_H4(135 	DOWNTO 128) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_CHUC(7 DOWNTO 0);
										 
	LCD_H4(143 	DOWNTO 136) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_DONVI(23 DOWNTO 16);
	LCD_H4(151 	DOWNTO 144) <= X"20" WHEN ENA_CP='0' ELSE  LCD_MA_DONVI(15 DOWNTO 8);
	LCD_H4(159 	DOWNTO 152) <= X"20" WHEN ENA_CP='0' ELSE LCD_MA_DONVI(7 DOWNTO 0);

end Behavioral;

