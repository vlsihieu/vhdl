
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY LCD_SOLON_TRAITIM IS 
	PORT ( CKHT : IN STD_LOGIC;
			 BTN_N: IN STD_LOGIC_VECTOR ( 1 DOWNTO 0);
			 LEDR: OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			 DS18B20: INOUT STD_LOGIC;
			 LCD_E: OUT STD_LOGIC;
			 LCD_RS: OUT STD_LOGIC;
			 LCD_RW: OUT STD_LOGIC;
			 LCD_ON: OUT STD_LOGIC;
			 LCD_BLON: OUT STD_LOGIC;			 
			 LCD_DB: OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0));
END LCD_SOLON_TRAITIM;
ARCHITECTURE PMH OF LCD_SOLON_TRAITIM IS 
--LCD 
SIGNAL LCD_HANG_1: STD_LOGIC_VECTOR ( 127 DOWNTO 0);
SIGNAL LCD_HANG_2: STD_LOGIC_VECTOR ( 127 DOWNTO 0);
signal DONVI,CHUC: std_logic_vector ( 3 downto 0);
SIGNAL DONVI_ND,CHUC_ND: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
SIGNAL LCD_MA_TO_CHUC,LCD_MA_TO_DONVI: STD_LOGIC_VECTOR ( 47 DOWNTO 0);
SIGNAL LCD_MA_TO_CHUC_ND,LCD_MA_TO_DONVI_ND: STD_LOGIC_VECTOR ( 47 DOWNTO 0);
--NHIET DO 
SIGNAL DS_PRESENT : STD_LOGIC;
SIGNAL NHIETDO: STD_LOGIC_VECTOR ( 7 DOWNTO 0);
SIGNAL TEMPERATURE : STD_LOGIC_VECTOR ( 11 DOWNTO 0);
-- NUT NHAN 
SIGNAL RST : STD_LOGIC;
SIGNAL MODE,MODE_CDLH: STD_LOGIC;
-- TIN HIEU
SIGNAL OE:STD_LOGIC_VECTOR ( 2 DOWNTO 0);
-- DEM
SIGNAL DEM: STD_LOGIC_VECTOR ( 7 DOWNTO 0 );
SIGNAL ENA_DB : STd_LOGIC;
BEGIN
	RST <= NOT BTN_N(0);
	MODE <= NOT BTN_N(1);
	NHIETDO <= TEMPERATURE (11 DOWNTO 4);
	LEDR( 3 DOWNTO 0) <= TEMPERATURE ( 3 DOWNTO 0);
   LCD_ON <= '1';
	LCD_RW <= '0';
CHIA_10ENA: ENTITY WORK.CHIA_10ENA	
	PORT MAP ( CKHT =>CKHT,
				  ENA2HZ=> ENA_DB);
DS18B20_TEMPERATURE : ENTITY WORK.DS18B20_TEMPERATURE -- DO NHIET DO 
	PORT MAP ( CKHT => CKHT,
					DS18B20 => DS18B20,
					RST => RST,
					DS_PRESENT => DS_PRESENT,
					TEMPERATURE_OUT => TEMPERATURE);
HEXTOBCD_ND: ENTITY WORK.HEXTOBCD_8BIT -- GIAI MA NHIET DO 
	PORT  MAP ( SOHEX8BIT => NHIETDO,
					DONVI => DONVI_ND,
					CHUC => CHUC_ND);
MACH_DEM: ENTITY WORK.DEM_8BIT -- DEM GH
	PORT MAP ( CKHT => CKHT,
				  ENA_DB => ENA_DB,
				  OE => OE,
				  RST => RST,
				  Q => DEM );
HEXTOBCD_DEM: ENTITY WORK.HEXTOBCD_8BIT -- GIAI MA DEM GIOI HAN 
	PORT MAP ( SOHEX8BIT => DEM,
				  DONVI => DONVI,
				  CHUC => CHUC);		
CD_LAM_HEP_BTN_MODE : ENTITY WORK.CD_LAM_HEP_BTN-- NUT NHAN MODE 
	PORT MAP ( CKHT => CKHT,
				  BTN => MODE,
				  BTN_CDLH => MODE_CDLH);
DIEUKHIEN_MODE: ENTITY WORK.DIEUKHIEN_MODE--DIEU KHIEN CHE DO OE 
	PORT MAP ( CKHT => CKHT,
				  MODE_CDLH => MODE_CDLH,
				  RST => RST,
				  OE => OE);
LCD_KHOITAO_HIENTHI: ENTITY WORK.LCD_KHOITAO_HIENTHI_CGRAM_SO_TO --
	PORT MAP (  LCD_DB => LCD_DB,
					LCD_RS => LCD_RS,
					LCD_E => LCD_E,
					LCD_RST => RST,
					LCD_CK => CKHT,
					OE => OE,
					LCD_HANG_1 => LCD_HANG_1,
					LCD_HANG_2 => LCD_HANG_2
	);
LCD_GAN_DULIEU_SO_TO: ENTITY WORK.LCD_GAN_DULIEU_3SO_TO--
	PORT MAP(	LCD_MA_TO_DONVI => LCD_MA_TO_DONVI,
					LCD_MA_TO_CHUC => LCD_MA_TO_CHUC,
					LCD_MA_TO_DONVI_ND => LCD_MA_TO_DONVI_ND,
					LCD_MA_TO_CHUC_ND => LCD_MA_TO_CHUC_ND,
					OE => OE,
					DONVI_ND=> DONVI_ND,
					CHUC_ND=> CHUC_ND,
					DONVI=> DONVI,
					CHUC=> CHUC,
					LCD_HANG_1 => LCD_HANG_1,
					LCD_HANG_2 => LCD_HANG_2
	);	  
LCD_GIAI_MA_DV_DEM: ENTITY WORK.LCD_GIAI_MA_DV
	PORT MAP ( DONVI_GM => DONVI,
				  CHUC_GM  => CHUC  ,
				  LCD_MA_TO_DONVI => LCD_MA_TO_DONVI,
				  LCD_MA_TO_CHUC => LCD_MA_TO_CHUC);
LCD_GIAI_MA_DV_ND: ENTITY WORK.LCD_GIAI_MA_DV
	PORT MAP ( DONVI_GM => DONVI_ND,
				  CHUC_GM  => CHUC_ND  ,
				  LCD_MA_TO_DONVI => LCD_MA_TO_DONVI_ND,
				  LCD_MA_TO_CHUC => LCD_MA_TO_CHUC_ND);
	END PMH;