library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
entity LCD_GAN_DULIEU_HIENTHI_NN is
    Port ( 	H1_9,H1_10,H1_12, H1_13, H1_15, H1_16, H1_7: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	
				GIATRI_MOD: IN STD_LOGIC_VECTOR(1 DOWNTO 0);
				NN: IN STD_LOGIC;
				LCD_HANG_1, LCD_HANG_2 : out  STD_LOGIC_VECTOR (127 downto 0));
end LCD_GAN_DULIEU_HIENTHI_NN;

architecture Behavioral of LCD_GAN_DULIEU_HIENTHI_NN is

begin
PROCESS(NN,GIATRI_MOD)
BEGin
IF(GIATRI_MOD="00") THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="01" AND NN='0') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="01" AND NN='1') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="10" AND NN='0') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="10" AND NN='1') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="11" AND NN='0') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
ELSIF (GIATRI_MOD="11" AND NN='1') THEN
	LCD_HANG_1(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('L'),8);
	LCD_HANG_1(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_1(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_1(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(':'),8);
	LCD_HANG_1(55 DOWNTO 48)	<= X"3" & H1_7;
	LCD_HANG_1(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(71 DOWNTO 64)	<= X"3" & H1_9;
	LCD_HANG_1(79 DOWNTO 72)	<= X"3" & H1_10;
	LCD_HANG_1(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(95 DOWNTO 88)	<= X"3" & H1_12;
	LCD_HANG_1(103 DOWNTO 96)	<= X"3" & H1_13;
	LCD_HANG_1(111 DOWNTO 104)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1(119 DOWNTO 112)	<= X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120)	<= X"3" & H1_16;
	
	LCD_HANG_2(7 DOWNTO 0)		<=	CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);
	LCD_HANG_2(15 DOWNTO 8)		<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('T'),8);
	LCD_HANG_2(23 DOWNTO 16)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('O'),8);
	LCD_HANG_2(31 DOWNTO 24)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_2(39 DOWNTO 32)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('N'),8);
	LCD_HANG_2(47 DOWNTO 40)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_2(55 DOWNTO 48)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('K'),8);
	LCD_HANG_2(63 DOWNTO 56)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(71 DOWNTO 64)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(79 DOWNTO 72)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(87 DOWNTO 80)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('4'),8);
	LCD_HANG_2(95 DOWNTO 88)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2(103 DOWNTO 96)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('3'),8);
	LCD_HANG_2(111 DOWNTO 104)<=  CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(119 DOWNTO 112)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('2'),8);
	LCD_HANG_2(127 DOWNTO 120)	<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('*'),8);	
END IF;
END PROCESS;
end Behavioral;