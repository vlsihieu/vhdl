LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;



ENTITY LED_STD_PST_A IS
PORT ( CKHT,RST,ENA_SS,ENA_DB,ON_PST,OFF_TSP:IN STD_LOGIC;
		Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END LED_STD_PST_A;

ARCHITECTURE THAN OF LED_STD_PST_A IS
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN Q_REG <= (OTHERS => '0');
	ELSIF FALLING_EDGE(CKHT) THEN Q_REG<=Q_NEXT;
	END IF;
END PROCESS;

PROCESS(ENA_DB,ON_PST,OFF_TSP,Q_REG,ENA_SS)
BEGIN
	Q_NEXT <= Q_REG;
	IF ENA_DB = '1' THEN
		IF ENA_SS = '1' THEN
			IF ON_PST = '1' THEN Q_NEXT <= Q_REG(6 DOWNTO 0) & NOT Q_REG(7);
			ELSIF OFF_TSP = '1' THEN Q_NEXT <= NOT Q_REG(0) & Q_REG(7 DOWNTO 1);
			END IF;
		ELSE
--			Q_NEXT <= (OTHERS => '0');
         Q_NEXT <= Q_REG;
		END IF;
	END IF;
END PROCESS;
	Q <= Q_REG;		
--Q <= Q_REG WHEN ENA_SS = '1' ELSE (OTHERS => '0');
END THAN;
