LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CD_4BTN IS
	PORT ( CKHT: IN STD_LOGIC;
			BTN_N: 	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			BTN0,BTN1,BTN2,BTN3: 	OUT STD_LOGIC
		   );
END CD_4BTN;

ARCHITECTURE BEHAVIOR OF CD_4BTN IS

BEGIN
CD_BTN_BTN0: ENTITY WORK.BTN
	PORT MAP(	CKHT 		=> CKHT,
					BTN 		=> NOT BTN_N(0),
					Q => BTN0
				);
CD_BTN_BTN1: ENTITY WORK.BTN
	PORT MAP(	CKHT 		=> CKHT,
					BTN 		=> NOT BTN_N(1),
					Q => BTN1
				);
CD_BTN_BTN2: ENTITY WORK.BTN
	PORT MAP(	CKHT 		=> CKHT,
					BTN 		=> NOT BTN_N(2),
					Q => BTN2
				);
CD_BTN_BTN3: ENTITY WORK.BTN
	PORT MAP(	CKHT 		=> CKHT,
					BTN 		=> NOT BTN_N(3),
					Q => BTN3
				);
				
					
	
	
	
	
END BEHAVIOR;