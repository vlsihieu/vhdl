library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;

entity LED_DSDC_TSP is
	Port ( CKHT,RST,ENA_DB,OE,CP: in STD_LOGIC;
			 Q: out STD_LOGIC_VECTOR(7 DOWNTO 0));
end LED_DSDC_TSP;
architecture Behavioral of LED_DSDC_TSP is
SIGNAL Q_REG,Q_NEXT: STD_LOGIC_VECTOR(7 DOWNTO 0);
begin
	PROCESS(CKHT,RST)
	BEGIN
		IF 	RST='1' 					THEN Q_REG <="10000000";
		ELSIF FALLING_EDGE(CKHT) 	THEN Q_REG <=Q_NEXT;
		END IF;
	END PROCESS;
	
	Q_NEXT <= "10000000" WHEN OE='0' AND CP = '0' ELSE
				 Q_REG(0) & Q_REG(7 DOWNTO 1)  WHEN ENA_DB ='1' AND OE='1' AND CP = '1' ELSE 
				 Q_REG;
				 
	Q <= Q_REG WHEN OE='1' AND CP = '1'  ELSE 
	    (OTHERS =>'0');
end Behavioral;