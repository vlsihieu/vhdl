library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity DEM_GIOPHUTGIAY is
    Port ( CKHT, RST, ENA_DB,ENA_UP, ENA_DW, ENA_CHINH : in  STD_LOGIC;
	 GT_MOD: STD_LOGIC_VECTOR(1 DOWNTO 0);
           GIAY, PHUT : out  STD_LOGIC_VECTOR (5 downto 0);
           GIO : out  STD_LOGIC_VECTOR (4 downto 0));
end DEM_GIOPHUTGIAY;

architecture Behavioral of DEM_GIOPHUTGIAY is
	SIGNAL GIAY_NEXT, GIAY_REG: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL PHUT_NEXT, PHUT_REG: STD_LOGIC_VECTOR(5 DOWNTO 0);
	SIGNAL GIO_NEXT, GIO_REG: STD_LOGIC_VECTOR(4 DOWNTO 0);
begin

	PROCESS(CKHT, RST)
	BEGIN
		IF RST='1' THEN 	GIAY_REG <= (OTHERS => '0');
								PHUT_REG <= (OTHERS => '0');
								GIO_REG  <= (OTHERS => '0');
		ELSIF FALLING_EDGE(CKHT) THEN GIAY_REG <= GIAY_NEXT;
											PHUT_REG <= PHUT_NEXT;
											GIO_REG  <= GIO_NEXT;
											
		END IF;
	END PROCESS;
	--===============================================
	PROCESS(GIAY_REG, ENA_DB,GT_MOD,ENA_UP,ENA_DW,ENA_CHINH)
	BEGIN
		GIAY_NEXT <= GIAY_REG;
		IF ENA_DB = '1' THEN
			IF GIAY_REG = "111011" THEN	GIAY_NEXT <= (OTHERS => '0');
			ELSE								GIAY_NEXT			<= GIAY_REG +1;
			END IF;
		ELSIF GT_MOD="01" AND ENA_UP='1' AND ENA_CHINH='1' THEN
			IF GIAY_REG = "111011" THEN	GIAY_NEXT <= (OTHERS => '0');
			ELSE								GIAY_NEXT			<= GIAY_REG +1;
			END IF;
		ELSIF GT_MOD="01" AND ENA_DW='1' AND ENA_CHINH='1' THEN
			IF GIAY_REG = "000000" THEN	GIAY_NEXT <=  "111011";
			ELSE								GIAY_NEXT			<= GIAY_REG -1;
			END IF;
			END IF;
	END PROCESS;
	--===============================================
	PROCESS(GIAY_REG, PHUT_REG,ENA_DB,GT_MOD,ENA_UP,ENA_DW,ENA_CHINH)
	BEGIN
		PHUT_NEXT <= PHUT_REG;
		IF ENA_DB = '1' AND GIAY_REG="111011" THEN
			IF PHUT_REG = "111011" THEN	PHUT_NEXT <= (OTHERS => '0');
			ELSE								PHUT_NEXT			<= PHUT_REG +1;
			END IF;
		ELSIF GT_MOD="10" AND ENA_UP='1' AND ENA_CHINH='1' THEN
			IF PHUT_REG = "111011" THEN	PHUT_NEXT <= (OTHERS => '0');
			ELSE								PHUT_NEXT			<= PHUT_REG +1;
			END IF;
		ELSIF GT_MOD="10" AND ENA_DW='1' AND ENA_CHINH='1' THEN
			IF PHUT_REG = "000000" THEN	PHUT_NEXT <= "111011";
			ELSE								PHUT_NEXT			<= PHUT_REG -1;
			END IF;
			END IF;
	END PROCESS;
	--=================================================
	PROCESS(GIAY_REG,GIO_REG, PHUT_REG,ENA_DB,GT_MOD,ENA_UP,ENA_DW,ENA_CHINH)
	BEGIN
		GIO_NEXT <= GIO_REG;
		IF ENA_DB = '1' AND GIAY_REG="111011" AND PHUT_REG = "111011" THEN
			IF GIO_REG = "10111" THEN	GIO_NEXT <= (OTHERS => '0');
			ELSE								GIO_NEXT			<= GIO_REG +1;
			END IF;
		ELSIF GT_MOD="11" AND ENA_UP='1' AND ENA_CHINH='1' THEN
			IF GIO_REG = "10111" THEN	GIO_NEXT <= (OTHERS => '0');
			ELSE								GIO_NEXT			<= GIO_REG +1;
			END IF;
		ELSIF GT_MOD="11" AND ENA_DW='1' AND ENA_CHINH='1' THEN
			IF GIO_REG = "00000" THEN	GIO_NEXT <= "10111";
			ELSE								GIO_NEXT			<= GIO_REG -1;
			END IF;
			END IF;
	END PROCESS;
	--=================================================
	GIAY	<= GIAY_REG;
	PHUT	<= PHUT_REG;
	GIO	<= GIO_REG;
end Behavioral;