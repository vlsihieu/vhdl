-- CHUONG TRINH CHIA XUNG CHO CAC BAI

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CHIA_10ENA IS 
	PORT( CKHT:   IN STD_LOGIC;
			ENA_UD : IN STD_LOGIC;
			ENA1KHZ : OUT STD_LOGIC;
			ENA_CK : OUT STD_LOGIC 
		  );
END CHIA_10ENA;
 
ARCHITECTURE BEHAVIORAL OF CHIA_10ENA IS

--SIGNAL ENA2HZ  : STD_LOGIC; 
SIGNAL ENA20HZ  : STD_LOGIC;  
SIGNAL ENA10HZ  : STD_LOGIC; 

CONSTANT N : INTEGER := 50000000;


SIGNAL D10HZ_REG,  D10HZ_NEXT   : INTEGER RANGE 0 TO N/10   := 1;
SIGNAL D20HZ_REG,  D20HZ_NEXT   : INTEGER RANGE 0 TO N/20   := 1;
SIGNAL D1KHZ_REG,  D1KHZ_NEXT   : INTEGER RANGE 0 TO N/1000 := 1;

BEGIN
-- OUTPUT LOGIC

	ENA1KHZ   <='1' WHEN D1KHZ_REG = N/(1000*2)  	  	ELSE '0';
	ENA20HZ   <='1' WHEN D20HZ_REG = N/(20*2)          ELSE '0';
	ENA10HZ   <='1' WHEN D10HZ_REG = N/(10*2)          ELSE '0';  

   ENA_CK    <= ENA20HZ WHEN ENA_UD = '1' ELSE
	             ENA10HZ;
	
-- REGISTER
PROCESS( CKHT)
BEGIN	
		IF FALLING_EDGE (CKHT) THEN D10HZ_REG   <= D10HZ_NEXT;
											 D20HZ_REG   <= D20HZ_NEXT;
											 D1KHZ_REG   <= D1KHZ_NEXT;

		END IF;
	END PROCESS;
	
-- NEXT STATE LOGIC

D10HZ_NEXT <= 1 WHEN D10HZ_REG = N/10 ELSE
						   D10HZ_REG +1;  

D20HZ_NEXT <= 1 WHEN D20HZ_REG = N/20 ELSE
						   D20HZ_REG +1;
--
D1KHZ_NEXT <= 1 WHEN D1KHZ_REG = N/1000 ELSE
						   D1KHZ_REG +1;

END BEHAVIORAL;
	