LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY DEM_2SO IS
PORT (CKHT,RST :IN STD_LOGIC;
		DONVI_A  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CHUC_A   :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DONVI_B  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CHUC_B   :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		ENA_DB   :IN STD_LOGIC;
		ENA_SS,ENA_UD   :IN STD_LOGIC;
		DONVI,CHUC      : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	   );
END DEM_2SO;

ARCHITECTURE THAN OF DEM_2SO IS
SIGNAL DONVI_REG, DONVI_NEXT : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG, CHUC_NEXT   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
BEGIN
PROCESS(CKHT,RST,DONVI_A,CHUC_A)
BEGIN
	IF RST='1'   THEN DONVI_REG <= DONVI_A;
							CHUC_REG  <= CHUC_A;
	ELSIF FALLING_EDGE(CKHT) THEN DONVI_REG  <= DONVI_NEXT;
											CHUC_REG   <= CHUC_NEXT;
	END IF;
END PROCESS;

PROCESS(DONVI_REG,CHUC_REG,ENA_SS,ENA_DB,ENA_UD,DONVI_A,DONVI_B,CHUC_A,CHUC_B)
BEGIN
-- KHI ENA_SS =0 DUNG CHUONG TRINH 
	DONVI_NEXT <= DONVI_REG;
	CHUC_NEXT  <= CHUC_REG;
--	DONVI_NEXT <= DONVI_A;
--	CHUC_NEXT  <= CHUC_A;
--------------------------
 IF ( CHUC_A >= CHUC_B) THEN  DONVI_NEXT <= DONVI_REG;
                                CHUC_NEXT <= CHUC_REG;
 ELSIF  (CHUC_A < CHUC_B) THEN
	IF (ENA_DB = '1' AND ENA_SS = '1' )THEN
	       
         IF (ENA_UD = '0' ) THEN 
				IF DONVI_REG = DONVI_B AND CHUC_REG = CHUC_B THEN DONVI_NEXT <= DONVI_A;
																				  CHUC_NEXT  <= CHUC_A;
				ELSIF DONVI_REG /= X"9" THEN DONVI_NEXT <= DONVI_REG + 1;
				ELSE							  
				   DONVI_NEXT <= X"0";
					IF CHUC_REG /= X"9" THEN CHUC_NEXT <= CHUC_REG + 1;
					ELSE							 CHUC_NEXT <= X"0";
					END IF;
				END IF;
			ELSE
				IF DONVI_REG = DONVI_A AND CHUC_REG = CHUC_A THEN DONVI_NEXT <= DONVI_B;
																				  CHUC_NEXT  <= CHUC_B;
				ELSIF DONVI_REG/= X"0" THEN DONVI_NEXT <= DONVI_REG - 1;
				ELSE 							 
				   DONVI_NEXT <= X"9";
					IF CHUC_REG /= X"0" THEN CHUC_NEXT <= CHUC_REG - 1;
					ELSE							 CHUC_NEXT <= X"9";
					END IF;
				END IF;
			END IF;   
	END IF;
 END IF;
END PROCESS;
					  
DONVI <= DONVI_REG ;
CHUC  <= CHUC_REG ;
	
END THAN;
