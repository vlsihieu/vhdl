LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY DIEUKHIEN_LED_3S IS 
	PORT ( Q_LED: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			 DEM : IN STD_LOGIC_VECTOR ( 5 DOWNTO 0);
			 NHIETDO: IN STD_LOGIC_VECTOR ( 7 DOWNTO 0);
			 LED : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0)
			 );
END DIEUKHIEN_LED_3S;
ARCHITECTURE PMH OF DIEUKHIEN_LED_3S IS 
SIGNAL Q: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
signal gt_dem : std_logic_vector(7 downto 0);
BEGIN
   gt_dem <= "00" & dem;
	PROCESS(gt_DEM,NHIETDO,Q_LED)
	BEGIN
		IF ( gt_DEM >= NHIETDO ) THEN Q <= Q_LED ;
		ELSIF ( gt_DEM = NHIETDO + "00001111") THEN Q <= "0000";
		END IF;
	END PROCESS;
	LED <= Q;
END PMH;		