
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity UART is
    Port ( CKHT : IN STD_LOGIC;
	        BTN0 : IN STD_LOGIC;
			  SW0  : IN STD_LOGIC;
			  UART_RX :  IN STD_LOGIC;
			  UART_TX : OUT STD_LOGIC;
			  LCD_E: OUT STD_LOGIC;
			  LCD_RS: OUT STD_LOGIC;
			  LCD_P: OUT STD_LOGIC;
			  LCD_DB: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
           SSEG : out  STD_LOGIC_VECTOR (7 downto 0);
           ANODE : out  STD_LOGIC_VECTOR (7 downto 0)
			  );
end UART;

architecture Behavioral of UART is
SIGNAL RST,ENA1KHZ  :  STD_LOGIC;
SIGNAL LCD_HANG_1_R : STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_HANG_1_N:  STD_LOGIC_VECTOR (159 downto 0);
--SIGNAL LCD_HANG_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

SIGNAL UART_TX_FULL : STD_LOGIC;
SIGNAL UART_RX_EMPTY: STD_LOGIC;

SIGNAL UART_RECV_DATA: STD_LOGIC_VECTOR (7 downto 0);
SIGNAL UART_TRANS_DATA: STD_LOGIC_VECTOR (7 downto 0);
SIGNAL UART_ENA_TX: STD_LOGIC;
SIGNAL UART_ENA_RD: STD_LOGIC;

SIGNAL ENA_DB: STD_LOGIC;
SIGNAL ENA_RX: STD_LOGIC;

SIGNAL DEM: STD_LOGIC_VECTOR (7 downto 0);
SIGNAL DONVI: STD_LOGIC_VECTOR (3 downto 0);
SIGNAL CHUC: STD_LOGIC_VECTOR (3 downto 0);
SIGNAL TRAM: STD_LOGIC_VECTOR (3 downto 0);

SIGNAL LCD_H2 : STD_LOGIC_VECTOR(159 DOWNTO 0);
SIGNAL DAU_CHAM_8LED:STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL ENA_GIAIMA_8LED:STD_LOGIC_VECTOR(7 DOWNTO 0);
begin
RST <= not BTN0;

ENA_RX <= CKHT;
LCD_P <='1';

DAU_CHAM_8LED		<=X"FF";    -- "11111111"
ENA_GIAIMA_8LED	<= "00000111";   ---"00000011" -- KHI THEM LED PHAI SUA LAI
	
IC1: ENTITY WORK.CHIA_10ENA
   PORT MAP(CKHT =>CKHT,
	         ENA10HZ => ENA_DB,
				ENA1KHZ => ENA1KHZ
				);

IC2: ENTITY WORK.UART_CONTROLLER
   PORT MAP(CKHT =>CKHT,
	         RST  => RST,
				UART_RX => UART_RX,
				UART_TX => UART_TX,
				FIFO_UART_RX_ENA_RD => UART_ENA_RD,
				FIFO_UART_RX_DATA_RD => UART_RECV_DATA,
				FIFO_UART_RX_EMPTY   => UART_RX_EMPTY,

				FIFO_UART_TX_ENA_WR => UART_ENA_TX,
				FIFO_UART_TX_DATA_WR => UART_TRANS_DATA,
				FIFO_UART_TX_FULL   => UART_TX_FULL
				);

--------------------				
PROCESS(UART_TX_FULL,ENA_DB,SW0,DEM)
BEGIN
  UART_TRANS_DATA <= DEM;
  IF UART_TX_FULL = '0' THEN
     UART_ENA_TX <= ENA_DB AND SW0; -- TAO XUNG PHAT
  ELSE
     UART_ENA_TX <='0';
  END IF;
END PROCESS;
----------------------
UART_ENA_RD <= ENA_RX AND ( NOT UART_RX_EMPTY);

PROCESS(CKHT,RST)
BEGIN
  IF RST = '1' THEN
     LCD_HANG_1_R <= X"2020202020202020202020202020202020202020";
  ELSIF FALLING_EDGE(CKHT) THEN LCD_HANG_1_R <= LCD_HANG_1_N;
  END IF;
END PROCESS;

LCD_HANG_1_N <=  UART_RECV_DATA & LCD_HANG_1_R(159 DOWNTO 8)
                 WHEN UART_ENA_RD = '1'
					  ELSE LCD_HANG_1_R;
------------------------
IC3: ENTITY WORK.DEM_8BIT
   PORT MAP(CKHT =>CKHT,
	         RST  => RST,
				ENA_SS => SW0,
	         ENA_DB => ENA_DB,
				DEM => DEM
				);
IC4 : ENTITY WORK.HEXTOBCD_8BIT
		PORT MAP(	SOHEX8BIT	=> DEM,
						DONVI			=> DONVI,
						CHUC			=> CHUC,
						TRAM 			=> TRAM);
						
IC5 : ENTITY WORK.LCD_20X4_GAN_DULIEU_3SO
		PORT MAP(	H2_17			=> TRAM,
						H2_18			=> CHUC,
						H2_19			=> DONVI,
						LCD_H2		=> LCD_H2
						);
						
IC6: ENTITY WORK.LCD_20X4_KHOITAO_HIENTHI
		PORT MAP(	LCD_DB	=> LCD_DB,
						LCD_RS	=> LCD_RS,
						LCD_E		=> LCD_E,
						LCD_RST	=> BTN0,
						LCD_CK	=> CKHT,
						LCD_H1	=> LCD_HANG_1_R,
						LCD_H2	=> LCD_H2
						);

HIENTHI_2LED: ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
		PORT MAP(CKHT => CKHT,
					ENA1KHZ => ENA1KHZ,
					LED70 => DONVI,
					LED71 => CHUC,
					LED72 => TRAM,
					LED73 => X"F",
					LED74 => X"F",
					LED75 => X"F",
					LED76 => X"F",
					LED77 => X"F",
					
					DC_8LED  => DAU_CHAM_8LED,
					ENA_8LED => ENA_GIAIMA_8LED,
					ANODE => ANODE,
					SSEG => SSEG);
end Behavioral;

