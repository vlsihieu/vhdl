LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DICH_LCD_BTN IS 
	PORT ( CKHT : IN STD_LOGIC;
			 BTN: IN STD_LOGIC_VECTOR ( 1 DOWNTO 0);
			 LCD_E: OUT STD_LOGIC;
			 LCD_RS: OUT STD_LOGIC;
			 LCD_RW: OUT STD_LOGIC;
			 LCD_DB: OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0)
			 );
END DICH_LCD_BTN;
ARCHITECTURE PMH OF DICH_LCD_BTN IS 
SIGNAL MODE,MODE_CDLH,RST: STD_LOGIC;
--
SIGNAL OE: STD_LOGIC;
SIGNAL LCD_HANG_1: STD_LOGIC_VECTOR ( 127 DOWNTO 0);
SIGNAL LCD_HANG_2: STD_LOGIC_VECTOR ( 127 DOWNTO 0);
BEGIN
	RST  <= NOT BTN(0);
	MODE <= NOT BTN(1);
--	LCD_ON <= '1';
	LCD_RW <= '0';
	OE <= '1' ;
IC0 : ENTITY WORK.CD_LAM_HEP_BTN--SS
	PORT MAP ( CKHT => CKHT,
				  BTN => MODE,
				  BTN_CDLH => MODE_CDLH
				  );
IC1: ENTITY WORK.LCD_GAN_DULIEU_3SO_TO--
	PORT MAP(	RST => RST,
					CKHT => CKHT,
					OE => OE,
					MODE_CDLH => MODE_CDLH,
					LCD_HANG_1 => LCD_HANG_1,
					LCD_HANG_2 =>LCD_HANG_2);
IC2: ENTITY WORK.LCD_KHOITAO_HIENTHI_CGRAM_SO_TO --
	PORT MAP ( LCD_DB => LCD_DB,
					LCD_RS => LCD_RS,
					LCD_E => LCD_E,
					LCD_RST => RST,
					LCD_CK => CKHT,
					LCD_HANG_1 => LCD_HANG_1,
					LCD_HANG_2 => LCD_HANG_2
	);
END PMH;