LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY BTVN_SO8 IS 
	PORT ( CKHT, BTN0 : IN STD_LOGIC;
			 LED : OUT STD_LOGIC_VECTOR ( 7 DOWNTO 0));
END BTVN_SO8;

ARCHITECTURE BEHAVIORAL OF BTVN_SO8 IS 
SIGNAL  RST: STD_LOGIC;
SIGNAL  ENA_DB: STD_LOGIC;
SIGNAL Q_SD_PST, Q_SD_TSP : STD_LOGIC_VECTOR  ( 7 DOWNTO 0 );
SIGNAL OE : STD_LOGIC_VECTOR( 1 DOWNTO 0 );
BEGIN 
	
	LED <= Q_SD_PST OR Q_SD_TSP;
	RST <= NOT BTN0 ;
				 
CHIA_10ENA : ENTITY WORK.CHIA_10ENA 
		PORT MAP ( CKHT => CKHT,
		           OE => OE,
						ENA_CK => ENA_DB);
						
LED_SANGDON_PST: ENTITY WORK.LED_SANGDON_PST 
		PORT MAP ( CKHT => CKHT,
						RST => RST,
						ENA_DB => ENA_DB,
						OE => OE(0),
						Q => Q_SD_PST);
						
LED_SANGDON_TSP: ENTITY WORK.LED_SANGDON_TSP
		PORT MAP ( CKHT => CKHT,
						RST => RST,
						ENA_DB => ENA_DB,
						OE => OE(1),
						Q => Q_SD_TSP);
						
						
DIEUKHIEN_CHOPHEP : ENTITY WORK.DIEUKHIEN_CHOPHEP
		PORT MAP (  CKHT => CKHT,
						RST => RST,
						ENA_DB=> ENA_DB,
						OE => OE);
	
END BEHAVIORAL;
