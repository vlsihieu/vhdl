LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DEM_2SO IS
PORT (CKHT,RST :IN STD_LOGIC;
		DONVI_A  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CHUC_A   :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		DONVI_B  :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		CHUC_B   :IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		ENA_DB   :IN STD_LOGIC;
		ena_ud   : in std_logic;
		ENA_SS,OE   :IN STD_LOGIC;
		DONVI,CHUC    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END DEM_2SO;

ARCHITECTURE THAN OF DEM_2SO IS
SIGNAL DONVI_REG, DONVI_NEXT : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG, CHUC_NEXT   : STD_LOGIC_VECTOR(3 DOWNTO 0);  
SIGNAL DONVI_REG_A, DONVI_NEXT_A : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_A, CHUC_NEXT_A   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
BEGIN
PROCESS(CKHT,RST,DONVI_A,CHUC_A)
BEGIN
	IF RST='1'  THEN
	  if (ena_ud = '1' ) then
	       donvi_reg <= donvi_a;
			 chuc_reg  <= chuc_a;
	  else
	       donvi_reg <= donvi_b;
			 chuc_reg  <= chuc_b;
	  end if;
	ELSIF FALLING_EDGE(CKHT) THEN DONVI_REG  <= DONVI_NEXT;
											CHUC_REG   <= CHUC_NEXT;
											DONVI_REG_A  <= DONVI_NEXT_A;
											CHUC_REG_A   <= CHUC_NEXT_A;
	END IF;
END PROCESS;

PROCESS(ena_ud,DONVI_REG,CHUC_REG,DONVI_REG_A,CHUC_REG_A,ENA_SS,ENA_DB,DONVI_A,DONVI_B,CHUC_A,CHUC_B,OE)
BEGIN
	DONVI_NEXT <= DONVI_REG;
	CHUC_NEXT  <= CHUC_REG;
	DONVI_NEXT_A <= DONVI_REG_A;
	CHUC_NEXT_A <= CHUC_REG_A;
	IF OE = '1' THEN 
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN
            if (ena_ud = '1' ) then			
					IF DONVI_REG_A = DONVI_B AND CHUC_REG_A = CHUC_B THEN DONVI_NEXT_A <= DONVI_A;
																					  CHUC_NEXT_A  <= CHUC_A;
					ELSIF DONVI_REG_A /= X"9" THEN DONVI_NEXT_A <= DONVI_REG_A + 1;
					ELSE							  DONVI_NEXT_A <= X"0";
						IF CHUC_REG_A /= X"9" THEN CHUC_NEXT_A <= CHUC_REG_A + 1;
						ELSE							 CHUC_NEXT_A <= X"0";
						END IF;
					END IF;
				 else
				   donvi_next_a <= donvi_reg_a;
					chuc_next_a <= chuc_reg_a;
				 end if;
			END IF;
		END IF;
	ELSE
	-- KHONG CHO PHEP THI HIEN THI 00 NHUNG KHI CHO PHEP THI DEM TU A
		DONVI_NEXT_A <= DONVI_A;
		CHUC_NEXT_A  <= CHUC_A;
		DONVI_NEXT <= X"0";
		CHUC_NEXT  <= X"0";
	END IF;
END PROCESS;
					  
	DONVI <= DONVI_REG_A WHEN OE = '1' ELSE
				DONVI_REG;
	CHUC  <= CHUC_REG_A WHEN  OE = '1' ELSE
				CHUC_REG;
END THAN;
