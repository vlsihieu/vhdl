LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIEUKHIEN_MODE IS
PORT (CKHT : IN STD_LOGIC;
      RST : IN STD_LOGIC;
--		ENA_DB : IN STD_LOGIC; 
		SW :IN STD_LOGIC;
		OE : OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END DIEUKHIEN_MODE;

ARCHITECTURE BEHAVIORAL OF DIEUKHIEN_MODE IS

SIGNAL DEM_N,DEM_R : INTEGER RANGE 0 TO 3 := 0 ;
BEGIN

PROCESS ( CKHT, RST)
	BEGIN 
		IF RST = '1'              THEN DEM_R <= 0;
		ELSIF FALLING_EDGE(CKHT ) THEN DEM_R <= DEM_N;
		END IF ;
END PROCESS;


DEM_N <= DEM_R + 1 WHEN SW = '1' AND DEM_R <3  ELSE	
			0 			 WHEN SW = '1' AND DEM_R =3 ELSE
			DEM_R ;

			
PROCESS (DEM_R,RST)
BEGIN
		OE<="000"; -- tung bit dai dien cho tung chuong trinh 0 1 2
   	IF(RST='1')     THEN OE<=  "000";           -- DE RESET
		ELSIF DEM_R = 0 THEN OE <= "000"; 	 -- DEM PST 
		ELSIF DEM_R = 1 THEN OE <= "001";   -- DEM TSP
		ELSIF DEM_R = 2 THEN OE <= "010";   -- DICH 1 LED
		ELSIF DEM_R = 3 THEN OE <= "100";   -- DICH 1 LED
		END IF;
		
END PROCESS;
END BEHAVIORAL;
