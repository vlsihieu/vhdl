library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.std_logic_unsigned.all;
USE IEEE.NUMERIC_STD.ALL;


entity DEM_3BIT_GIAIMA is
    Port ( CKHT,RST,ENA : in  STD_LOGIC;
           OE : out  STD_LOGIC_VECTOR (3 downto 0));
end DEM_3BIT_GIAIMA;

architecture Behavioral of DEM_3BIT_GIAIMA is
SIGNAL Q_REG,Q_NEXT : STD_LOGIC_VECTOR( 2 DOWNTO 0);
begin
   PROCESS(CKHT, RST)
	BEGIN
	  IF RST='1' THEN Q_REG <= (OTHERS =>'0');
	  ELSIF FALLING_EDGE (CKHT) THEN Q_REG <= Q_NEXT;
	  END IF;
	END PROCESS;
  Q_NEXT <= Q_REG + 1 WHEN ENA ='1' ELSE
				"000"     WHEN Q_REG = "101" ELSE 
            Q_REG;
  PROCESS(Q_REG,RST)
  BEGIN
		OE<="0000";
		IF RST='1' THEN OE <="0000";
		ELSIF Q_REG="000" THEN OE <="0000";
		ELSIF Q_REG="001" THEN OE <="0001";
		ELSIF Q_REG="010" THEN OE <="0010";
		ELSIF Q_REG="011" THEN OE <="0100";
		ELSIF Q_REG="100" THEN OE <="1000";
		END IF;
	END PROCESS;
end Behavioral;

