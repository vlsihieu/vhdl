LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_5BIT IS
	PORT (CKHT : IN STD_LOGIC;
	      RST : IN STD_LOGIC;
			ENA_SS : IN STD_LOGIC;
			ENA_DB: IN STD_LOGIC;
			Q: OUT STD_LOGIC_VECTOR(4 DOWNTO 0)
			);
END DEM_5BIT;

ARCHITECTURE A OF DEM_5BIT IS
SIGNAL Q_REG : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
SIGNAL Q_NEXT: STD_LOGIC_VECTOR(4 DOWNTO 0);
BEGIN
---------------------
	PROCESS (CKHT, RST)
	BEGIN
		IF RST='1' 				     THEN Q_REG <= "01011";
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG<= Q_NEXT;
		END IF;
	END PROCESS;
-------------------------	
	Q_NEXT <= "01011" WHEN (Q_REG = "11111") AND ENA_SS = '1' AND ENA_DB = '1' ELSE 
				 Q_REG + 1 WHEN ENA_DB='1' AND ENA_SS = '1' ELSE 
				 Q_REG;
--------------------------				 
	Q <= Q_REG;
END A;