LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DIEUKHIEN_SS IS 
	PORT ( CKHT : in std_logic;
	       ENA_DB: IN STD_LOGIC;
			 Q: OUT STD_LOGIC
			 );
END DIEUKHIEN_SS;
ARCHITECTURE PMH OF DIEUKHIEN_SS IS 
SIGNAL DEM_REG, DEM_NEXT:  STD_LOGIC;
BEGIN
	--REGISTER 
	PROCESS(CKHT)
	BEGIN
		IF FALLING_EDGE (CKHT) THEN DEM_REG <= DEM_NEXT ;
		END IF ;
	END PROCESS;
 -- NEXT STATE 
	DEM_NEXT <= NOT DEM_REG WHEN ENA_DB ='1' ELSE 
						 DEM_REG;
	Q <= DEM_REG;
END PMH;
