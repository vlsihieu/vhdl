LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
---- vi no co 4 lua chon  ---> oe 2bit
ENTITY DIEUKHIEN_MODE IS
	PORT (CKHT,RST,MODE_CDLH: IN STD_LOGIC;
			OE: OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
		   );
END DIEUKHIEN_MODE;

ARCHITECTURE A OF DIEUKHIEN_MODE IS
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(1 DOWNTO 0):="00";
BEGIN
	PROCESS (CKHT, RST)
	BEGIN
		IF RST='1' 				     THEN Q_REG <= (OTHERS =>'0');
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG<= Q_NEXT;
		END IF;
	END PROCESS;
	
	Q_NEXT <= Q_REG +1 WHEN MODE_CDLH='1' ELSE 
				 Q_REG;		 
	OE <= Q_REG;
END A;