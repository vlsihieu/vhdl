-- CHUONG TRINH CHIA XUNG CHO CAC BAI

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY CHIA_10ENA IS 
	PORT( CKHT:   IN STD_LOGIC;
			ENA_UD : IN STD_LOGIC;
			ENA1KHZ : OUT STD_LOGIC;
			ENA_CK : OUT STD_LOGIC 
		  );
END CHIA_10ENA;
 
ARCHITECTURE BEHAVIORAL OF CHIA_10ENA IS

--SIGNAL ENA2HZ  : STD_LOGIC; 
SIGNAL ENA2HZ  : STD_LOGIC;  
SIGNAL ENA5HZ  : STD_LOGIC; 

CONSTANT N : INTEGER := 50000000;


SIGNAL D2HZ_REG,  D2HZ_NEXT   : INTEGER RANGE 0 TO N/2   := 1;
SIGNAL D5HZ_REG,  D5HZ_NEXT   : INTEGER RANGE 0 TO N/5   := 1;
SIGNAL D1KHZ_REG,  D1KHZ_NEXT   : INTEGER RANGE 0 TO N/1000 := 1;

BEGIN
-- OUTPUT LOGIC

	ENA1KHZ   <='1' WHEN D1KHZ_REG = N/(1000*2)  	  	ELSE '0';
	ENA5HZ   <='1' WHEN D5HZ_REG = N/(5*2)          ELSE '0';
	ENA2HZ   <='1' WHEN D2HZ_REG = N/(2*2)          ELSE '0';  

   ENA_CK    <= ENA2HZ WHEN ENA_UD = '1' ELSE
	             ENA5HZ;
	
-- REGISTER
PROCESS( CKHT)
BEGIN	
		IF FALLING_EDGE (CKHT) THEN D5HZ_REG   <= D5HZ_NEXT;
											 D2HZ_REG   <= D2HZ_NEXT;
											 D1KHZ_REG   <= D1KHZ_NEXT;

		END IF;
	END PROCESS;
	
-- NEXT STATE LOGIC

D2HZ_NEXT <= 1 WHEN D2HZ_REG = N/2 ELSE
						   D2HZ_REG +1;  

D5HZ_NEXT <= 1 WHEN D5HZ_REG = N/5 ELSE
						   D5HZ_REG +1;
--
D1KHZ_NEXT <= 1 WHEN D1KHZ_REG = N/1000 ELSE
						   D1KHZ_REG +1;

END BEHAVIORAL;
	