LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DEM_2SO IS
PORT (CKHT,RST :IN STD_LOGIC;
		OE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
		ENA_DB   :IN STD_LOGIC;
		ENA_SS   :IN STD_LOGIC;
		DONVI,CHUC    : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END DEM_2SO;

ARCHITECTURE THAN OF DEM_2SO IS
SIGNAL DONVI_REG, DONVI_NEXT : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG, CHUC_NEXT   : STD_LOGIC_VECTOR(3 DOWNTO 0);  
SIGNAL DONVI_REG_0, DONVI_NEXT_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_0, CHUC_NEXT_0   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL DONVI_REG_1, DONVI_NEXT_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_1, CHUC_NEXT_1   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL DONVI_REG_2, DONVI_NEXT_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_2, CHUC_NEXT_2   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL DONVI_REG_3, DONVI_NEXT_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_3, CHUC_NEXT_3   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL DONVI_REG_4, DONVI_NEXT_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_4, CHUC_NEXT_4   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
SIGNAL DONVI_REG_5, DONVI_NEXT_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG_5, CHUC_NEXT_5   : STD_LOGIC_VECTOR(3 DOWNTO 0); 
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN DONVI_REG <= (OTHERS => '0');
							CHUC_REG  <= (OTHERS => '0');
	ELSIF FALLING_EDGE(CKHT) THEN DONVI_REG  <= DONVI_NEXT;
											CHUC_REG   <= CHUC_NEXT;
											DONVI_REG_0  <= DONVI_NEXT_0;
											CHUC_REG_0   <= CHUC_NEXT_0;
											DONVI_REG_1  <= DONVI_NEXT_1;
											CHUC_REG_1   <= CHUC_NEXT_1;
											DONVI_REG_2  <= DONVI_NEXT_2;
											CHUC_REG_2   <= CHUC_NEXT_2;
											DONVI_REG_3  <= DONVI_NEXT_3;
											CHUC_REG_3   <= CHUC_NEXT_3;
											DONVI_REG_4  <= DONVI_NEXT_4;
											CHUC_REG_4   <= CHUC_NEXT_4;
											DONVI_REG_5  <= DONVI_NEXT_5;
											CHUC_REG_5   <= CHUC_NEXT_5;
	END IF;
END PROCESS;

PROCESS(DONVI_REG,CHUC_REG,ENA_SS,ENA_DB,OE,DONVI_REG_0,CHUC_REG_0,DONVI_REG_1,CHUC_REG_1,DONVI_REG_2,CHUC_REG_2,DONVI_REG_3,CHUC_REG_3,DONVI_REG_4,CHUC_REG_4,DONVI_REG_5,CHUC_REG_5)
BEGIN
	DONVI_NEXT <= DONVI_REG;
	CHUC_NEXT  <= CHUC_REG;
	DONVI_NEXT_0 <= DONVI_REG_0;
	CHUC_NEXT_0  <= CHUC_REG_0;
	DONVI_NEXT_1 <= DONVI_REG_1;
	CHUC_NEXT_1  <= CHUC_REG_1;
	DONVI_NEXT_2 <= DONVI_REG_2;
	CHUC_NEXT_2  <= CHUC_REG_2;
	DONVI_NEXT_3 <= DONVI_REG_3;
	CHUC_NEXT_3  <= CHUC_REG_3;
	DONVI_NEXT_4 <= DONVI_REG_4;
	CHUC_NEXT_4  <= CHUC_REG_4;
	DONVI_NEXT_5 <= DONVI_REG_5;
	CHUC_NEXT_5  <= CHUC_REG_5;
	
	IF OE(0) = '1' THEN
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_0 = X"0" AND CHUC_REG_0 = X"2" THEN DONVI_NEXT_0 <= DONVI_REG_0;
																			    CHUC_NEXT_0  <= CHUC_REG_0;
				ELSIF DONVI_REG_0 /= X"9" THEN DONVI_NEXT_0 <= DONVI_REG_0 + 1;
				ELSE							  DONVI_NEXT_0 <= X"0";
					IF CHUC_REG_0 /= X"9" THEN CHUC_NEXT_0 <= CHUC_REG_0 + 1;
					ELSE							 CHUC_NEXT_0 <= X"0";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSIF OE(1) = '1' THEN 
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_1 = X"0" AND CHUC_REG_1 = X"4" THEN DONVI_NEXT_1 <= DONVI_REG_1;
																			CHUC_NEXT_1  <= CHUC_REG_1;
				ELSIF DONVI_REG_1 /= X"9" THEN DONVI_NEXT_1 <= DONVI_REG_1 + 1;
				ELSE							  DONVI_NEXT_1 <= X"0";
					IF CHUC_REG_1 /= X"9" THEN CHUC_NEXT_1 <= CHUC_REG_1 + 1;
					ELSE							 CHUC_NEXT_1 <= X"0";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSIF OE(2) = '1' THEN
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_2 = X"1" AND CHUC_REG_2 = X"1" THEN DONVI_NEXT_2 <= DONVI_REG_2;
																			CHUC_NEXT_2  <= CHUC_REG_2;
				ELSIF DONVI_REG_2 /= X"0" THEN DONVI_NEXT_2 <= DONVI_REG_2 - 1;
				ELSE							  DONVI_NEXT_2 <= X"9";
					IF CHUC_REG_2 /= X"0" THEN CHUC_NEXT_2 <= CHUC_REG_2 - 1;
					ELSE							 CHUC_NEXT_2 <= X"9";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSIF OE(3) = '1' THEN
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_3 = X"0" AND CHUC_REG_3 = X"0" THEN DONVI_NEXT_3 <= DONVI_REG_3;
																			CHUC_NEXT_3  <= CHUC_REG_3;
				ELSIF DONVI_REG_3 /= X"0" THEN DONVI_NEXT_3 <= DONVI_REG_3 - 1;
				ELSE							  DONVI_NEXT_3 <= X"9";
					IF CHUC_REG_3 /= X"0" THEN CHUC_NEXT_3 <= CHUC_REG_3 - 1;
					ELSE							 CHUC_NEXT_3 <= X"9";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSIF OE(4) = '1' THEN	
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_4 = X"0" AND CHUC_REG_4 = X"6" THEN DONVI_NEXT_4 <= DONVI_REG_4;
																			CHUC_NEXT_4  <= CHUC_REG_4;
				ELSIF DONVI_REG_4 /= X"8" THEN DONVI_NEXT_4 <= DONVI_REG_4 + 2;
				ELSE							  DONVI_NEXT_4 <= X"0";
					IF CHUC_REG_4 /= X"6" THEN CHUC_NEXT_4 <= CHUC_REG_4 + 1;
					ELSE							 CHUC_NEXT_4 <= X"0";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSIF OE(5) = '1' THEN
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		IF ENA_DB = '1' THEN	
			IF ENA_SS = '1' THEN 
				IF DONVI_REG_5 = X"1" AND CHUC_REG_5 = X"0" THEN DONVI_NEXT_5 <= DONVI_REG_5;
																			CHUC_NEXT_5  <= CHUC_REG_5;
				ELSIF DONVI_REG_5 /= X"1" THEN DONVI_NEXT_5 <= DONVI_REG_5 - 2;
				ELSE							  DONVI_NEXT_5 <= X"9";
					IF CHUC_REG_5 /= X"0" THEN CHUC_NEXT_5 <= CHUC_REG_5 - 1;
					ELSE							 CHUC_NEXT_5 <= X"9";
					END IF;
				END IF;
			END IF;
		END IF;
	ELSE 
		DONVI_NEXT <= X"0";
		CHUC_NEXT <= X"0";
		DONVI_NEXT_0 <= X"0";
		CHUC_NEXT_0  <= X"0";
		DONVI_NEXT_1 <= X"1";
		CHUC_NEXT_1  <= X"2";
		DONVI_NEXT_2 <= X"0";
		CHUC_NEXT_2  <= X"4";
		DONVI_NEXT_3 <= X"0";
		CHUC_NEXT_3  <= X"1";
		DONVI_NEXT_4 <= X"0";
		CHUC_NEXT_4  <= X"0";
		DONVI_NEXT_5 <= X"9";
		CHUC_NEXT_5  <= X"5";
	END IF;
END PROCESS;
	

		
	DONVI <= DONVI_REG_0 WHEN OE(0) = '1' ELSE
				DONVI_REG_1 WHEN OE(1) = '1' ELSE
				DONVI_REG_2 WHEN OE(2) = '1' ELSE
				DONVI_REG_3 WHEN OE(3) = '1' ELSE
				DONVI_REG_4 WHEN OE(4) = '1' ELSE
				DONVI_REG_5 WHEN OE(5) = '1' ELSE
				DONVI_REG;
	CHUC  <= CHUC_REG_0 WHEN OE(0) = '1' ELSE
				CHUC_REG_1 WHEN OE(1) = '1' ELSE
				CHUC_REG_2 WHEN OE(2) = '1' ELSE
				CHUC_REG_3 WHEN OE(3) = '1' ELSE
				CHUC_REG_4 WHEN OE(4) = '1' ELSE
				CHUC_REG_5 WHEN OE(5) = '1' ELSE
				CHUC_REG;
	
END THAN;
