LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DEM_2SO IS
PORT (CKHT,RST   :IN STD_LOGIC;
		ENA_DB     :IN STD_LOGIC;
		ENA_SS     :IN STD_LOGIC;
		ENA_UP     :IN STD_LOGIC;
		ENA_DW     :IN STD_LOGIC;
		DONVI,CHUC : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
	   );
END DEM_2SO;

ARCHITECTURE THAN OF DEM_2SO IS
SIGNAL DONVI_REG, DONVI_NEXT : STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC_REG, CHUC_NEXT   : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN DONVI_REG <= (OTHERS => '0');
							CHUC_REG  <= (OTHERS => '0');
	ELSIF FALLING_EDGE(CKHT) THEN DONVI_REG  <= DONVI_NEXT;
						 					CHUC_REG   <= CHUC_NEXT;
	END IF;
END PROCESS;

PROCESS(DONVI_REG,CHUC_REG,ENA_UP,ENA_DW,ENA_DB,ENA_SS)
BEGIN
	DONVI_NEXT <= DONVI_REG;
	CHUC_NEXT  <= CHUC_REG;
	IF ENA_SS = '1' THEN
		IF ENA_DB = '1' THEN	
			IF ENA_UP = '1' THEN 
					IF DONVI_REG = X"0" AND CHUC_REG = X"2" THEN DONVI_NEXT <= DONVI_REG;
																			   CHUC_NEXT  <= CHUC_REG;
					ELSIF DONVI_REG /= X"9" THEN DONVI_NEXT <= DONVI_REG + 1;
					ELSE							  
					   DONVI_NEXT <= X"0";
						IF CHUC_REG /= X"9" THEN CHUC_NEXT <= CHUC_REG + 1;
						ELSE							 CHUC_NEXT <= X"0";
						END IF;
					END IF;
			ELSIF ENA_DW = '1' THEN
					IF DONVI_REG = X"0" AND CHUC_REG = X"0" THEN DONVI_NEXT <= DONVI_REG;
																			   CHUC_NEXT  <= CHUC_REG;
					ELSIF DONVI_REG /= X"0" THEN DONVI_NEXT <= DONVI_REG - 1;
					ELSE							  
					   DONVI_NEXT <= X"9";
						IF CHUC_REG /= X"0" THEN CHUC_NEXT <= CHUC_REG - 1;
						ELSE							 CHUC_NEXT <= X"9";
						END IF;
					END IF;
			END IF;
		END IF;
	END IF;
END PROCESS;
					  
	DONVI <= DONVI_REG;
	CHUC  <= CHUC_REG;
	
END THAN;
