library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity LED_STD_PST is
    Port (CKHT, RST, OE, ENA_DB:   in      STD_LOGIC;
    		Q:      out     STD_LOGIC_VECTOR (5 downto 0));
end LED_STD_PST;

architecture Behavioral of LED_STD_PST is
SIGNAL 	Q_REG, Q_NEXT: STD_LOGIC_VECTOR(5 DOWNTO 0);
Begin
   PROCESS (CKHT, RST)
   BEGIN   
		IF  RST='1'             THEN    Q_REG	<=	(OTHERS => '0'); 
      ELSIF   FALLING_EDGE (CKHT)   THEN    Q_REG	<=	Q_NEXT;	
		END IF;
	END PROCESS;
	
	Q_NEXT <= Q_REG(4 DOWNTO 0) & NOT Q_REG(5) WHEN ENA_DB = '1' ELSE
				 Q_REG;
       
	Q <= Q_REG WHEN OE = '1' ELSE (OTHERS => '0'); 
end Behavioral;