LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DEM_GH_UD_2BTN IS
	PORT( CKHT, RST, UP : IN STD_LOGIC;
			DONVI_GH, CHUC_GH: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END DEM_GH_UD_2BTN;
ARCHITECTURE BEHAVIORAL OF DEM_GH_UD_2BTN IS
SIGNAL DONVI_REG, DONVI_NEXT, CHUC_REG, CHUC_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
--REGISTER
	PROCESS(CKHT, RST)
	BEGIN
		IF RST = '1' THEN DONVI_REG <= x"2";
								CHUC_REG <= x"0";
		ELSIF FALLING_EDGE(CKHT) THEN DONVI_REG <= DONVI_NEXT;
												CHUC_REG <= CHUC_NEXT;
		END IF;
	END PROCESS;
--NEXT STATE LOGIC
	PROCESS(DONVI_REG, CHUC_REG, UP)
	BEGIN
		DONVI_NEXT <= DONVI_REG;
		CHUC_NEXT  <= CHUC_REG;
			IF UP = '1' THEN
				IF CHUC_REG&DONVI_REG = X"82" THEN DONVI_NEXT <= X"2"; CHUC_NEXT <= X"0";
				ELSE
				   
				--IF DONVI_REG /= X"9" THEN DONVI_NEXT <= DONVI_REG + 20;
					--ELSE							  DONVI_NEXT <= X"0";
						IF CHUC_REG /= X"9" THEN CHUC_NEXT <= CHUC_REG +2;
						ELSE							 CHUC_NEXT <= X"0";
					END IF;
					END IF;
				
			END IF;
	END PROCESS;
--OUTPUT LOGIC
	DONVI_GH <= DONVI_REG;
	CHUC_GH <= CHUC_REG;
END BEHAVIORAL;