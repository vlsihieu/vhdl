LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY LCD_GAN_DULIEU_3SO_TO IS
	PORT(	H1_0,H1_1,H1_15,H1_16: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			H2_0,H2_1: IN STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			LCD_HANG_1: OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
			LCD_HANG_2: OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
			ENA_DB_TMP,CKHT,RST : IN STD_LOGIC;
			OE : IN STD_LOGIC_VECTOR ( 1 DOWNTO 0);
			CK2HZ: IN STD_LOGIC
	);
END LCD_GAN_DULIEU_3SO_TO;

ARCHITECTURE BEHAVIORAL OF LCD_GAN_DULIEU_3SO_TO IS
SIGNAL LCD_HANG_1_1: STD_LOGIC_VECTOR ( 239 DOWNTO 0);
SIGNAL LCD_HANG_1_1_TMP: STD_LOGIC_VECTOR ( 79 DOWNTO 0);
SIGNAL I_REG,I_NEXT : INTEGER RANGE 0 TO 256 := 0;
SIGNAL LCD_HANG_2_1,LCD_HANG_2_1_TMP: STD_LOGIC_VECTOR ( 127 DOWNTO 0);
BEGIN
	-- HANG1
	LCD_HANG_1(7 DOWNTO 0) <= X"3" & H1_0; --TT
	LCD_HANG_1(15 DOWNTO 8) <=X"3" & H1_1;--TT
	LCD_HANG_1(23 DOWNTO 16)<= X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0  WHEN OE="01" ELSE 
										X"3" & H1_1  WHEN OE="10" ELSE 
										X"3" & H1_0 ;
	LCD_HANG_1(31 DOWNTO 24) <=X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0 WHEN OE="01" ELSE 
										X"3" & H1_1 WHEN OE="10" ELSE 
										X"3" & H1_0 ;
	LCD_HANG_1(39 DOWNTO 32)<= X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0 WHEN OE="01" ELSE 
										X"3" & H1_1 WHEN OE="10" ELSE 
										X"3" & H1_0 ;
	--- CON PHAN DICH CHU MACH DEM BCD
	LCD_HANG_1(111 DOWNTO 88) <= X"202020"; -- DAU CACH 
	LCD_HANG_1(119 DOWNTO 112) <=X"3" & H1_15;
	LCD_HANG_1(127 DOWNTO 120) <=X"3" & H1_16;
	---------BIEN LCD_HANG_11
	LCD_HANG_1_1(7 DOWNTO 0) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(15 DOWNTO 8) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(23 DOWNTO 16) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(31 DOWNTO 24) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(39 DOWNTO 32) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(47 DOWNTO 40) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(55 DOWNTO 48) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(63 DOWNTO 56) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(71 DOWNTO 64) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_1_1(79 DOWNTO 72) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
   LCD_HANG_1_1(87 DOWNTO 80)  <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8);
	LCD_HANG_1_1(95 DOWNTO 88)  <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('A'),8);
	LCD_HANG_1_1(103 DOWNTO 96) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1_1(111 DOWNTO 104)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('H'),8);
	LCD_HANG_1_1(119 DOWNTO 112)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_HANG_1_1(127 DOWNTO 120)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('E'),8);
	LCD_HANG_1_1(135 DOWNTO 128) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('M'),8);
	LCD_HANG_1_1(143 DOWNTO 136) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('B'),8);
	LCD_HANG_1_1(151 DOWNTO 144) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('C'),8);
	LCD_HANG_1_1(159 DOWNTO 152) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('D'),8);
	LCD_HANG_1_1(167 DOWNTO 160) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(175 DOWNTO 168) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(183 DOWNTO 176) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(191 DOWNTO 184) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(199 DOWNTO 192) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(207 DOWNTO 200) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(215 DOWNTO 208) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(223 DOWNTO 216) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8); --
			LCD_HANG_1_1(231 DOWNTO 224) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
			LCD_HANG_1_1(239 DOWNTO 232) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	--- XU LY DICH HANG 1 ----------
	PROCESS(RST,CKHT)
	BEGIN
		IF (RST = '1' ) THEN I_REG <= 0;
		ELSIF FALLING_EDGE(CKHT) THEN I_REG <= I_NEXT;
		END IF;
	END PROCESS;
	I_NEXT <= 	0 WHEN I_REG = 160 AND ENA_DB_TMP = '1'  ELSE -- OE TAC DONG VAO DE DEM 
					I_REG + 8 WHEN ENA_DB_TMP = '1' ELSE
					I_REG;
	LCD_HANG_1_1_TMP <= LCD_HANG_1_1((I_REG+79) DOWNTO I_REG );
	------ HIEN THI HANG 1 ------------
	LCD_HANG_1(87 DOWNTO 40) <= LCD_HANG_1_1_TMP ( 47 DOWNTO 0);
	-- HANG2
	--------------------------HANG 2 ---------------------------
	LCD_HANG_2 ( 7 DOWNTO 0) <= X"3" & H2_0;
	LCD_HANG_2(15 DOWNTO 8) <= X"3" & H2_1;
	LCD_HANG_2(23 DOWNTO 16)<= X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0 WHEN OE="01" ELSE 
										X"3" & H1_1 WHEN OE="10" ELSE 
										X"3" & H1_0;
	LCD_HANG_2(31 DOWNTO 24)<= X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0 WHEN OE="01" ELSE 
										X"3" & H1_1 WHEN OE="10" ELSE 
										X"3" & H1_0 ;
	LCD_HANG_2(39 DOWNTO 32)<= X"3" & H2_1  WHEN OE="00" ELSE  -- XXX
										X"3" & H2_0 WHEN OE="01" ELSE 
										X"3" & H1_1 WHEN OE="10" ELSE 
										X"3" & H1_0 ;
	---- HIEN THI CHOP TAT HANG 2 
	LCD_HANG_2_1(7 DOWNTO 0) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(15 DOWNTO 8) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(23 DOWNTO 16) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(31 DOWNTO 24) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(39 DOWNTO 32) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(47 DOWNTO 40) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(55 DOWNTO 48) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(63 DOWNTO 56) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2_1(71 DOWNTO 64) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2_1(79 DOWNTO 72) <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('6'),8);
   LCD_HANG_2_1(87 DOWNTO 80)  <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2_1(95 DOWNTO 88)  <=CONV_STD_LOGIC_VECTOR(CHARACTER'POS('1'),8);
	LCD_HANG_2_1(103 DOWNTO 96) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('9'),8);
	LCD_HANG_2_1(111 DOWNTO 104)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('0'),8);
	LCD_HANG_2_1(119 DOWNTO 112)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('8'),8);
	LCD_HANG_2_1(127 DOWNTO 120)<= CONV_STD_LOGIC_VECTOR(CHARACTER'POS('7'),8);
	---- LCD__ HANG 2 
	LCD_HANG_2 ( 103 DOWNTO 40) <= LCD_HANG_2_1(63 DOWNTO 0) WHEN CK2HZ='1' ELSE 
											LCD_HANG_2_1(127 DOWNTO 64);
	LCD_HANG_2(111 DOWNTO 104) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(119 DOWNTO 112) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	LCD_HANG_2(127 DOWNTO 120) <= CONV_STD_LOGIC_VECTOR(CHARACTER'POS(' '),8);
	 -- MUON SANG VI TRI NAO THI CHO NO BANG X"00"
END BEHAVIORAL;
