LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY BTVN_SO7 IS
	PORT (CKHT : IN STD_LOGIC;
	      BTN  : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			LED : OUT STD_LOGIC_VECTOR( 7 DOWNTO 0));
END BTVN_SO7;

ARCHITECTURE BEHAVIORAL OF BTVN_SO7 IS
SIGNAL ENA_DB: STD_LOGIC ;
SIGNAL RST : STD_LOGIC;
SIGNAL BTN_N1 : STD_LOGIC;
SIGNAL ENA_TT : STD_LOGIC;
SIGNAL BTN_CDLH : STD_LOGIC;
SIGNAL BTN_MODE : STD_LOGIC;
SIGNAL Q_STD_PST : STD_LOGIC_VECTOR ( 7 DOWNTO 0);
SIGNAL Q_STD_TSP : STD_LOGIC_VECTOR ( 3 DOWNTO 0);
SIGNAL OE : STD_LOGIC_VECTOR( 1 DOWNTO 0 );

BEGIN 
	RST <=  NOT  BTN(0);
	BTN_MODE <= NOT BTN(1);

-- dem_1bit_btn
IC0 : ENTITY WORK.CD_LAM_HEP_BTN
		PORT  MAP ( CKHT => CKHT,
						BTN  =>  BTN_MODE, -- NGO VAO BTN CHUYEN CHE DO
						BTN_CDLH => BTN_CDLH);

IC1 : ENTITY WORK.DEM_1BIT
     PORT MAP ( CKHT => CKHT,
	             RST  => RST,
					 ENA_DB => BTN_CDLH,
					 Q     => ENA_TT );
            	  

IC2 : ENTITY WORK.CHIA_10ENA 
	PORT  MAP ( CKHT  => CKHT,
					ENA5HZ => ENA_DB);
			
IC3 : ENTITY WORK.LED_STD_PST 
	PORT MAP ( CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					OE => OE(0),
					Q => Q_STD_PST);
					
IC4 : ENTITY WORK.LED_STD_4LED_TSP 
	PORT MAP ( CKHT => CKHT,
					RST => RST,
					ENA_DB => ENA_DB,
					OE => OE(1),
					Q => Q_STD_TSP);
					
LED (5 DOWNTO 2) <=  Q_STD_PST(5 DOWNTO 2) OR Q_STD_TSP(3 DOWNTO 0);
LED (1 DOWNTO 0) <=  Q_STD_PST(1 DOWNTO 0);  
LED (7 DOWNTO 6) <=  Q_STD_PST(7 DOWNTO 6);
 OE <= "01" WHEN ENA_TT = '0' ELSE
		   "10" ;
					
					
END BEHAVIORAL;
