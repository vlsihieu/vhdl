LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY DEM_6BIT IS
	PORT (CKHT: IN STD_LOGIC;
	      RST : IN STD_LOGIC;
			ENA_DB: IN STD_LOGIC;
	      ENA_SS : IN STD_LOGIC;
			ena : out std_logic;
			Q: OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
		   );
END DEM_6BIT;

ARCHITECTURE A OF DEM_6BIT IS
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(5 DOWNTO 0);
BEGIN
	PROCESS (CKHT, RST)
	BEGIN
		IF RST='1' 				     THEN Q_REG <= (OTHERS =>'0');
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG<= Q_NEXT;
		END IF;
	END PROCESS;
	
	Q_NEXT <= "000000" WHEN Q_REG="110010" AND ENA_DB = '1' and ena_ss = '1' ELSE 
				 Q_REG +1 WHEN ENA_DB='1' and ena_ss = '1' ELSE 
				 Q_REG;					 
	Q <= Q_REG;
	ena <= '1' when (Q_REG = "110010") else
	       '0';
END A;