LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY xu_ly_choptat IS
      PORT (CKHT : IN STD_LOGIC;
		      ENA_DB : IN STD_LOGIC;
				ENA_SS: IN STD_LOGIC;
		      Q : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
				);
END xu_ly_choptat;
ARCHITECTURE PMH OF xu_ly_choptat IS
SIGNAL Q_REG : STD_LOGIC_VECTOR(3 DOWNTO 0):="0000";
signal Q_NEXT: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
 PROCESS(CKHT)
        BEGIN
				 IF FALLING_EDGE(CKHT) THEN Q_REG <= Q_NEXT;
				 END IF;
		  END PROCESS;
   Q_NEXT <= (OTHERS =>'0') WHEN ENA_SS='0' ELSE
              NOT(Q_REG)    WHEN ENA_SS='1' AND ENA_DB = '1' ELSE
				  Q_REG;
   Q <= Q_REG ;
END PMH; 