library ieee;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
ENTITY DIEUKHIEN_GH IS 
	PORT ( GT_MOD: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			 RST: IN STD_LOGIC;
			 ENA_UP: IN STD_LOGIC;
			 CKHT: IN STD_LOGIC;
			 GH_DV_TREN : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			 GH_DV_DUOI: OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			 GH_CHUC_TREN :  OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0);
			 GH_CHUC_DUOI : OUT STD_LOGIC_VECTOR ( 3 DOWNTO 0)
			);
END DIEUKHIEN_GH;
ARCHITECTURE PMH OF DIEUKHIEN_GH IS 
SIGNAL Q_REG1,Q_NEXT1: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
SIGNAL Q_REG2,Q_NEXT2: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
SIGNAL Q_REG3,Q_NEXT3: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
SIGNAL Q_REG4,Q_NEXT4: STD_LOGIC_VECTOR ( 3 DOWNTO 0);
BEGIN
	PROCESS (CKHT, RST)
	BEGIN
		IF RST='1' 				     THEN Q_REG1 <= (OTHERS =>'0');
												 Q_REG2 <= (OTHERS =>'0');
												 Q_REG3 <= (OTHERS =>'0');
												 Q_REG4 <= (OTHERS =>'0');											  
		ELSIF FALLING_EDGE (CKHT) THEN Q_REG1<= Q_NEXT1;
												 Q_REG2<= Q_NEXT2;
												 Q_REG3<= Q_NEXT3;
												 Q_REG4<= Q_NEXT4;
		END IF;
	END PROCESS;
	PROCESS(GT_MOD,ENA_UP,Q_REG1,Q_REG2,Q_REG3,Q_REG4)
	BEGIN
		Q_NEXT1 <= Q_REG1;
		Q_NEXT2 <= Q_REG2;
		Q_NEXT3 <= Q_REG3;
		Q_NEXT4 <= Q_REG4;
		IF GT_MOD="00" AND ENA_UP='1' THEN 
			IF Q_REG1="1001" THEN Q_NEXT1 <= "0000";
			ELSE Q_NEXT1 <= Q_REG1 + 1 ;
			END IF;
		ELSIF GT_MOD="01" AND ENA_UP='1' THEN 
			IF Q_REG2="1001" THEN Q_NEXT2 <= "0000";
			ELSE Q_NEXT2 <= Q_REG2 + 1 ;
			END IF;
		ELSIF GT_MOD="10" AND ENA_UP='1' THEN 
			IF Q_REG3="1001" THEN Q_NEXT3 <= "0000";
			ELSE Q_NEXT3 <= Q_REG3 + 1 ;
			END IF;
		ELSIF GT_MOD="11" AND ENA_UP='1' THEN 
			IF Q_REG4="1001" THEN Q_NEXT4 <= "0000";
			ELSE Q_NEXT4 <= Q_REG4 + 1 ;
			END IF;
		END IF;
	END PROCESS;
--	GH_DV_DUOI <= Q_REG1;
--	GH_CHUC_DUOI <= Q_REG2;
--	GH_DV_TREN <= Q_REG3;
--	GH_CHUC_TREN <= Q_REG4;
	GH_CHUC_TREN  <= Q_REG1;
	GH_DV_TREN <= Q_REG2;
	GH_CHUC_DUOI <= Q_REG3;
	GH_DV_DUOI <= Q_REG4;
END PMH;