LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DIEUKHIEN_CHOPHEP IS
PORT (CKHT,RST,ENA_DB :IN STD_LOGIC;
		OE : OUT STD_LOGIC_VECTOR(1 DOWNTO 0));
END DIEUKHIEN_CHOPHEP;

ARCHITECTURE BEHAVIORAL OF DIEUKHIEN_CHOPHEP IS
SIGNAL DEM_REG, DEM_NEXT: INTEGER RANGE 0 TO 73 := 0;
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN DEM_REG <= 0;
	ELSIF FALLING_EDGE(CKHT) THEN DEM_REG<=DEM_NEXT;
	END IF;
END PROCESS;

DEM_NEXT <= 0         WHEN DEM_REG = 73  AND ENA_DB ='1'   ELSE
			   DEM_REG+1 WHEN ENA_DB = '1'  ELSE
				DEM_REG;
				
PROCESS (DEM_REG,RST)
BEGIN
		OE<="00";
		IF(RST='1') THEN OE<="00";           -- DE RESET
		ELSIF DEM_REG <37 THEN OE <= "01"; 	 -- DEM PST 
		ELSE                    OE <= "10";   -- DEM TSP
		END IF;
END PROCESS;
END BEHAVIORAL;
