LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;



ENTITY LED_STD_PST_7 IS
PORT ( CKHT : IN STD_LOGIC;
       RST : IN STD_LOGIC;
		 ENA_DB  :IN STD_LOGIC;
		 ON_PST : IN STD_LOGIC;
		 OFF_TSP: IN STD_LOGIC;
		 OE : IN STD_LOGIC;
		 Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END LED_STD_PST_7;

ARCHITECTURE THAN OF LED_STD_PST_7 IS
SIGNAL Q_REG, Q_NEXT: STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
PROCESS(CKHT,RST)
BEGIN
	IF RST='1'   THEN Q_REG <= (OTHERS => '0');
	ELSIF FALLING_EDGE(CKHT) THEN Q_REG<=Q_NEXT;
	END IF;
END PROCESS;

PROCESS(ENA_DB,ON_PST,OFF_TSP,Q_REG,OE)
BEGIN
	Q_NEXT <= Q_REG;
	IF ENA_DB = '1' THEN
	  IF OE = '1' THEN 
		 IF ON_PST = '1' THEN 
		    IF (Q_REG = "11111111" ) THEN Q_NEXT <= Q_REG;
			 ELSE                         Q_NEXT <= Q_REG(6 DOWNTO 0) & NOT Q_REG(7);
			 END IF;
		 ELSIF OFF_TSP = '1' THEN 
		    IF (Q_REG = "00000000") THEN Q_NEXT <= Q_REG;
			 ELSE                         Q_NEXT <= NOT Q_REG(0) & Q_REG(7 DOWNTO 1);
			 END IF;
		 END IF;
	  END IF;
	END IF;
END PROCESS;
	Q <= Q_REG;		
--Q <= Q_REG WHEN ENA_SS = '1' ELSE (OTHERS => '0');
END THAN;
