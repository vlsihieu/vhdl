
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity CLOCK_DS18B20_LCD20X4_SO_TO_NHO is
    Port ( CKHT : in  STD_LOGIC;
           SW0 : in  STD_LOGIC;
			  BTN: in std_logic_vector(1 downto 0);
           LCD_P,LCD_E,LCD_RS : out  STD_LOGIC;
			  LCD_DB : out  STD_LOGIC_VECTOR (7 downto 0);
			  DS18B20 : INOUT STD_LOGIC;
			  LED : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
           ANODE : out  STD_LOGIC_VECTOR (7 downto 0);
           SSEG : out  STD_LOGIC_VECTOR (7 downto 0));
end CLOCK_DS18B20_LCD20X4_SO_TO_NHO;

architecture Behavioral of CLOCK_DS18B20_LCD20X4_SO_TO_NHO is
--DONGHO
SIGNAL LCD_H1:	STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_H2:	STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_H3:	STD_LOGIC_VECTOR (159 downto 0);
SIGNAL LCD_H4:	STD_LOGIC_VECTOR (159 downto 0);

SIGNAL LCD_MA_DV_GIO: STD_LOGIC_VECTOR(47 DOWNTO 0);

SIGNAL LCD_MA_CH_GIO: STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL GIAY, PHUT, GIO: STD_LOGIC_VECTOR(5 DOWNTO 0);
SIGNAL GIO5:				STD_LOGIC_VECTOR(4 DOWNTO 0);

SIGNAL CH_GIO, DV_GIO:	STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CH_PHUT, DV_PHUT:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL Ch_GIAY, DV_GIAY:STD_LOGIC_VECTOR(3 DOWNTO 0);
--NHIETDO
SIGNAL LCD_MA_DONVI: STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL LCD_MA_CHUC: 	STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL LCD_MA_TRAM: 	STD_LOGIC_VECTOR(47 DOWNTO 0);
SIGNAL DONVI:			STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL CHUC:			STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL TRAM:			STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LED0: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LED1: STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL LED2: STD_LOGIC_VECTOR(3 DOWNTO 0);

SIGNAL NHIETDO: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL GH_CHUC,GH_TRAM,GH_DONVI: STD_LOGIC_VECTOR( 3 DOWNTO 0);
SIGNAL DS_PRESENT: STD_LOGIC;
SIGNAL TEMPERATURE:  STD_LOGIC_VECTOR(11 DOWNTO 0);
SIGNAL ENA_DB,ENA_CK,ENA_CP,RST,ENA1KHZ: STD_LOGIC;
SIGNAL ND_GH: STD_LOGIC_VECTOR(7 DOWNTO 0);
--7SEG
SIGNAL 	DAU_CHAM_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL 	ENA_GIAIMA_8LED: STD_LOGIC_VECTOR(7 DOWNTO 0);
SIGNAL   OE: STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL   Q_STD_TNV,Q_STD_TTR: STD_LOGIC_VECTOR(15 DOWNTO 0);
begin

LCD_P	<= '1';
RST<=BTN(0);
GIO	<= '0'&GIO5;

NHIETDO	 <= TEMPERATURE(11 DOWNTO 4); 
ENA_CP <= '1' WHEN NHIETDO >= ND_GH ELSE '0';

DAU_CHAM_8LED	<=	X"FF";
ENA_GIAIMA_8LED	<= "11000000";
LED <= Q_STD_TNV OR Q_STD_TTR;	
	
OE<="01" WHEN ENA_CP='0' ELSE "10";
		
IC1: ENTITY WORK.LED_STD_TNV
PORT MAP( CKHT		=>CKHT,
			 RST		=>RST,
			 ENA_DB	=>  ENA_DB,
			 OE		=>OE(0),
			 Q			=>Q_STD_TNV);
			 
IC2: ENTITY WORK.LED_STD_TTR
PORT MAP( CKHT		=>CKHT,
			 RST		=>RST,
			 ENA_DB	=>  ENA_DB,
			 OE		=>OE(1),
			 Q			=>Q_STD_TTR);
			 
IC3: ENTITY WORK.DEBOUNCE_BTN
	PORT MAP (	CKHT		=> CKHT,
					BTN		=> BTN(1),
					DB_TICK	=> ENA_CK);
					
IC4: ENTITY WORK.DEM_8BIT
		PORT MAP( CKHT => CKHT,
					 RST => RST,
					 ENA_CK => ENA_CK,
					 ENA_DB=>ENA_DB,
					 Q => ND_GH);
					 
IC5: ENTITY WORK.HEXTOBCD_8BIT
	PORT MAP(	SOHEX8BIT	=> ND_GH,
					DONVI			=> GH_DONVI,
					CHUC			=> GH_CHUC,
					TRAM			=> GH_TRAM);
					
IC6:	ENTITY WORK.GIAIMA_HIENTHI_8LED_7DOAN
			PORT MAP (	CKHT				=>	CKHT,
							ENA1KHZ 			=> ENA1KHZ,
							LED70				=>	X"F",
							LED71				=>	X"F",
							LED72				=>	X"F",
							LED73				=>	X"F",
							LED74				=>	X"F",
							LED75				=>	X"F",
							LED76				=>	GH_DONVI,
							LED77				=>	GH_CHUC,							
							DAU_CHAM_8LED	=>	DAU_CHAM_8LED,							
							ENA_GIAIMA_8LED =>	ENA_GIAIMA_8LED,
							ANODE	=>	ANODE,
							SSEG	=>	SSEG);	
							
IC7: ENTITY WORK.DS18B20_TEMPERATURE
	PORT MAP(	CKHT			=> CKHT,
					RST			=> RST,
					DS18B20		=> DS18B20,
					DS_PRESENT	=> DS_PRESENT,
					TEMPERATURE	=> TEMPERATURE);
					
	PROCESS(DS_PRESENT, DONVI, CHUC, TRAM)
	BEGIN
		IF	(DS_PRESENT = '0') THEN		LED0	<= DONVI;
												LED1	<= CHUC;
												LED2  <= TRAM;
												
		ELSE					   			LED0	<= X"E";
												LED1	<= X"E";
												LED2	<= X"E";
		END IF;
	END PROCESS;
	
					
IC8: ENTITY WORK.HEXTOBCD_8BIT
	PORT MAP(	SOHEX8BIT	=> NHIETDO,
					DONVI			=> DONVI,
					CHUC			=> CHUC,
					TRAM			=> TRAM);
					
--------------NHIET DO --------------------					
IC9: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(	SO_GMA	=> LED0,
					LCD_MA_TO=> LCD_MA_DONVI);

IC10: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(	SO_GMA	=> LED1,
					LCD_MA_TO=> LCD_MA_CHUC);
--------------------------------------------
					
IC11: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(	SO_GMA	=> LED2,
					LCD_MA_TO=> LCD_MA_TRAM);	
					
IC12: ENTITY WORK.CHIA_10ENA
	PORT MAP(	CKHT		=> CKHT,
					ENA1KHZ	=>ENA1KHZ,
					ENA5HZ	=> ENA_DB);
					
IC13: ENTITY WORK.DEM_GIOPHUTGIAY
	PORT MAP(	CKHT		=> CKHT,
					RST		=> RST,
					ENA_DB	=> ENA_DB,
					GIO		=> GIO5,
					PHUT		=> PHUT,
					GIAY		=> GIAY);
					
IC14: ENTITY WORK.HEXTOBCD_6BIT
	PORT MAP(	SOHEX6BIT	=> GIO,
					DONVI			=> DV_GIO,
					CHUC			=> CH_GIO);
					
IC15: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(	SO_GMA	=> DV_GIO,
					LCD_MA_TO=> LCD_MA_DV_GIO);

IC16: ENTITY WORK.LCD_GIAI_MA_SO_TO
	PORT MAP(	SO_GMA	=> CH_GIO,
					LCD_MA_TO=> LCD_MA_CH_GIO);
					
					
IC17: ENTITY WORK.HEXTOBCD_6BIT
	PORT MAP(	SOHEX6BIT	=> PHUT,
					DONVI			=> DV_PHUT,
					CHUC			=> CH_PHUT);
					
IC18: ENTITY WORK.HEXTOBCD_6BIT
	PORT MAP(	SOHEX6BIT	=> GIAY,
					DONVI			=> DV_GIAY,
					CHUC			=> CH_GIAY);
					
IC19: ENTITY WORK.LCD_20X4_GAN_DULIEU_1SO_TO
	PORT MAP(	LCD_MA_DONVI	=> LCD_MA_DONVI,
					LCD_MA_CHUC		=> LCD_MA_CHUC,
					LCD_MA_TRAM		=> LCD_MA_TRAM,
					
					LCD_MA_CH_GIO		=> LCD_MA_CH_GIO,
					LCD_MA_DV_GIO		=> LCD_MA_DV_GIO,
					
					ENA_CP			   =>ENA_CP,
					ENA_TN				=>SW0,
					
					ND_TRAM			=>LED2,
					ND_CHUC			=>LED1,
					ND_DV				=>LED0,
					
					H1_12		=> CH_GIO,
					H1_13		=> DV_GIO,
					H1_15		=> CH_PHUT,
					H1_16		=> DV_PHUT,
					H1_18		=> CH_GIAY,
					H1_19		=> DV_GIAY,
					
					LCD_H1	=> LCD_H1,
					LCD_H2	=> LCD_H2,
					LCD_H3	=> LCD_H3,
					LCD_H4	=> LCD_H4);
					
IC20: ENTITY WORK.LCD_20X4_KHOITAO_HIENTHI_SO_TO
PORT MAP(	LCD_DB => LCD_DB,
				LCD_RS => LCD_RS,
				LCD_E => LCD_E,
				LCD_RST => RST,
				LCD_CK => CKHT,
				LCD_H1 => LCD_H1,
				LCD_H2 => LCD_H2,
				LCD_H3 => LCD_H3,
				LCD_H4 => LCD_H4);
				
end Behavioral;

